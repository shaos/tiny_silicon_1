magic
tech gf180mcuC
magscale 1 5
timestamp 1669961268
<< obsm1 >>
rect 40672 52767 149312 133497
<< metal2 >>
rect 5796 299760 5908 300480
rect 16884 299760 16996 300480
rect 27972 299760 28084 300480
rect 39060 299760 39172 300480
rect 50148 299760 50260 300480
rect 61236 299760 61348 300480
rect 72324 299760 72436 300480
rect 83412 299760 83524 300480
rect 94500 299760 94612 300480
rect 105588 299760 105700 300480
rect 116676 299760 116788 300480
rect 127764 299760 127876 300480
rect 138852 299760 138964 300480
rect 149940 299760 150052 300480
rect 161028 299760 161140 300480
rect 172116 299760 172228 300480
rect 183204 299760 183316 300480
rect 194292 299760 194404 300480
rect 205380 299760 205492 300480
rect 216468 299760 216580 300480
rect 227556 299760 227668 300480
rect 238644 299760 238756 300480
rect 249732 299760 249844 300480
rect 260820 299760 260932 300480
rect 271908 299760 272020 300480
rect 282996 299760 283108 300480
rect 294084 299760 294196 300480
rect 6636 -480 6748 240
rect 7588 -480 7700 240
rect 8540 -480 8652 240
rect 9492 -480 9604 240
rect 10444 -480 10556 240
rect 11396 -480 11508 240
rect 12348 -480 12460 240
rect 13300 -480 13412 240
rect 14252 -480 14364 240
rect 15204 -480 15316 240
rect 16156 -480 16268 240
rect 17108 -480 17220 240
rect 18060 -480 18172 240
rect 19012 -480 19124 240
rect 19964 -480 20076 240
rect 20916 -480 21028 240
rect 21868 -480 21980 240
rect 22820 -480 22932 240
rect 23772 -480 23884 240
rect 24724 -480 24836 240
rect 25676 -480 25788 240
rect 26628 -480 26740 240
rect 27580 -480 27692 240
rect 28532 -480 28644 240
rect 29484 -480 29596 240
rect 30436 -480 30548 240
rect 31388 -480 31500 240
rect 32340 -480 32452 240
rect 33292 -480 33404 240
rect 34244 -480 34356 240
rect 35196 -480 35308 240
rect 36148 -480 36260 240
rect 37100 -480 37212 240
rect 38052 -480 38164 240
rect 39004 -480 39116 240
rect 39956 -480 40068 240
rect 40908 -480 41020 240
rect 41860 -480 41972 240
rect 42812 -480 42924 240
rect 43764 -480 43876 240
rect 44716 -480 44828 240
rect 45668 -480 45780 240
rect 46620 -480 46732 240
rect 47572 -480 47684 240
rect 48524 -480 48636 240
rect 49476 -480 49588 240
rect 50428 -480 50540 240
rect 51380 -480 51492 240
rect 52332 -480 52444 240
rect 53284 -480 53396 240
rect 54236 -480 54348 240
rect 55188 -480 55300 240
rect 56140 -480 56252 240
rect 57092 -480 57204 240
rect 58044 -480 58156 240
rect 58996 -480 59108 240
rect 59948 -480 60060 240
rect 60900 -480 61012 240
rect 61852 -480 61964 240
rect 62804 -480 62916 240
rect 63756 -480 63868 240
rect 64708 -480 64820 240
rect 65660 -480 65772 240
rect 66612 -480 66724 240
rect 67564 -480 67676 240
rect 68516 -480 68628 240
rect 69468 -480 69580 240
rect 70420 -480 70532 240
rect 71372 -480 71484 240
rect 72324 -480 72436 240
rect 73276 -480 73388 240
rect 74228 -480 74340 240
rect 75180 -480 75292 240
rect 76132 -480 76244 240
rect 77084 -480 77196 240
rect 78036 -480 78148 240
rect 78988 -480 79100 240
rect 79940 -480 80052 240
rect 80892 -480 81004 240
rect 81844 -480 81956 240
rect 82796 -480 82908 240
rect 83748 -480 83860 240
rect 84700 -480 84812 240
rect 85652 -480 85764 240
rect 86604 -480 86716 240
rect 87556 -480 87668 240
rect 88508 -480 88620 240
rect 89460 -480 89572 240
rect 90412 -480 90524 240
rect 91364 -480 91476 240
rect 92316 -480 92428 240
rect 93268 -480 93380 240
rect 94220 -480 94332 240
rect 95172 -480 95284 240
rect 96124 -480 96236 240
rect 97076 -480 97188 240
rect 98028 -480 98140 240
rect 98980 -480 99092 240
rect 99932 -480 100044 240
rect 100884 -480 100996 240
rect 101836 -480 101948 240
rect 102788 -480 102900 240
rect 103740 -480 103852 240
rect 104692 -480 104804 240
rect 105644 -480 105756 240
rect 106596 -480 106708 240
rect 107548 -480 107660 240
rect 108500 -480 108612 240
rect 109452 -480 109564 240
rect 110404 -480 110516 240
rect 111356 -480 111468 240
rect 112308 -480 112420 240
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115164 -480 115276 240
rect 116116 -480 116228 240
rect 117068 -480 117180 240
rect 118020 -480 118132 240
rect 118972 -480 119084 240
rect 119924 -480 120036 240
rect 120876 -480 120988 240
rect 121828 -480 121940 240
rect 122780 -480 122892 240
rect 123732 -480 123844 240
rect 124684 -480 124796 240
rect 125636 -480 125748 240
rect 126588 -480 126700 240
rect 127540 -480 127652 240
rect 128492 -480 128604 240
rect 129444 -480 129556 240
rect 130396 -480 130508 240
rect 131348 -480 131460 240
rect 132300 -480 132412 240
rect 133252 -480 133364 240
rect 134204 -480 134316 240
rect 135156 -480 135268 240
rect 136108 -480 136220 240
rect 137060 -480 137172 240
rect 138012 -480 138124 240
rect 138964 -480 139076 240
rect 139916 -480 140028 240
rect 140868 -480 140980 240
rect 141820 -480 141932 240
rect 142772 -480 142884 240
rect 143724 -480 143836 240
rect 144676 -480 144788 240
rect 145628 -480 145740 240
rect 146580 -480 146692 240
rect 147532 -480 147644 240
rect 148484 -480 148596 240
rect 149436 -480 149548 240
rect 150388 -480 150500 240
rect 151340 -480 151452 240
rect 152292 -480 152404 240
rect 153244 -480 153356 240
rect 154196 -480 154308 240
rect 155148 -480 155260 240
rect 156100 -480 156212 240
rect 157052 -480 157164 240
rect 158004 -480 158116 240
rect 158956 -480 159068 240
rect 159908 -480 160020 240
rect 160860 -480 160972 240
rect 161812 -480 161924 240
rect 162764 -480 162876 240
rect 163716 -480 163828 240
rect 164668 -480 164780 240
rect 165620 -480 165732 240
rect 166572 -480 166684 240
rect 167524 -480 167636 240
rect 168476 -480 168588 240
rect 169428 -480 169540 240
rect 170380 -480 170492 240
rect 171332 -480 171444 240
rect 172284 -480 172396 240
rect 173236 -480 173348 240
rect 174188 -480 174300 240
rect 175140 -480 175252 240
rect 176092 -480 176204 240
rect 177044 -480 177156 240
rect 177996 -480 178108 240
rect 178948 -480 179060 240
rect 179900 -480 180012 240
rect 180852 -480 180964 240
rect 181804 -480 181916 240
rect 182756 -480 182868 240
rect 183708 -480 183820 240
rect 184660 -480 184772 240
rect 185612 -480 185724 240
rect 186564 -480 186676 240
rect 187516 -480 187628 240
rect 188468 -480 188580 240
rect 189420 -480 189532 240
rect 190372 -480 190484 240
rect 191324 -480 191436 240
rect 192276 -480 192388 240
rect 193228 -480 193340 240
rect 194180 -480 194292 240
rect 195132 -480 195244 240
rect 196084 -480 196196 240
rect 197036 -480 197148 240
rect 197988 -480 198100 240
rect 198940 -480 199052 240
rect 199892 -480 200004 240
rect 200844 -480 200956 240
rect 201796 -480 201908 240
rect 202748 -480 202860 240
rect 203700 -480 203812 240
rect 204652 -480 204764 240
rect 205604 -480 205716 240
rect 206556 -480 206668 240
rect 207508 -480 207620 240
rect 208460 -480 208572 240
rect 209412 -480 209524 240
rect 210364 -480 210476 240
rect 211316 -480 211428 240
rect 212268 -480 212380 240
rect 213220 -480 213332 240
rect 214172 -480 214284 240
rect 215124 -480 215236 240
rect 216076 -480 216188 240
rect 217028 -480 217140 240
rect 217980 -480 218092 240
rect 218932 -480 219044 240
rect 219884 -480 219996 240
rect 220836 -480 220948 240
rect 221788 -480 221900 240
rect 222740 -480 222852 240
rect 223692 -480 223804 240
rect 224644 -480 224756 240
rect 225596 -480 225708 240
rect 226548 -480 226660 240
rect 227500 -480 227612 240
rect 228452 -480 228564 240
rect 229404 -480 229516 240
rect 230356 -480 230468 240
rect 231308 -480 231420 240
rect 232260 -480 232372 240
rect 233212 -480 233324 240
rect 234164 -480 234276 240
rect 235116 -480 235228 240
rect 236068 -480 236180 240
rect 237020 -480 237132 240
rect 237972 -480 238084 240
rect 238924 -480 239036 240
rect 239876 -480 239988 240
rect 240828 -480 240940 240
rect 241780 -480 241892 240
rect 242732 -480 242844 240
rect 243684 -480 243796 240
rect 244636 -480 244748 240
rect 245588 -480 245700 240
rect 246540 -480 246652 240
rect 247492 -480 247604 240
rect 248444 -480 248556 240
rect 249396 -480 249508 240
rect 250348 -480 250460 240
rect 251300 -480 251412 240
rect 252252 -480 252364 240
rect 253204 -480 253316 240
rect 254156 -480 254268 240
rect 255108 -480 255220 240
rect 256060 -480 256172 240
rect 257012 -480 257124 240
rect 257964 -480 258076 240
rect 258916 -480 259028 240
rect 259868 -480 259980 240
rect 260820 -480 260932 240
rect 261772 -480 261884 240
rect 262724 -480 262836 240
rect 263676 -480 263788 240
rect 264628 -480 264740 240
rect 265580 -480 265692 240
rect 266532 -480 266644 240
rect 267484 -480 267596 240
rect 268436 -480 268548 240
rect 269388 -480 269500 240
rect 270340 -480 270452 240
rect 271292 -480 271404 240
rect 272244 -480 272356 240
rect 273196 -480 273308 240
rect 274148 -480 274260 240
rect 275100 -480 275212 240
rect 276052 -480 276164 240
rect 277004 -480 277116 240
rect 277956 -480 278068 240
rect 278908 -480 279020 240
rect 279860 -480 279972 240
rect 280812 -480 280924 240
rect 281764 -480 281876 240
rect 282716 -480 282828 240
rect 283668 -480 283780 240
rect 284620 -480 284732 240
rect 285572 -480 285684 240
rect 286524 -480 286636 240
rect 287476 -480 287588 240
rect 288428 -480 288540 240
rect 289380 -480 289492 240
rect 290332 -480 290444 240
rect 291284 -480 291396 240
rect 292236 -480 292348 240
rect 293188 -480 293300 240
<< obsm2 >>
rect 1246 299730 5766 299810
rect 5938 299730 16854 299810
rect 17026 299730 27942 299810
rect 28114 299730 39030 299810
rect 39202 299730 50118 299810
rect 50290 299730 61206 299810
rect 61378 299730 72294 299810
rect 72466 299730 83382 299810
rect 83554 299730 94470 299810
rect 94642 299730 105558 299810
rect 105730 299730 116646 299810
rect 116818 299730 127734 299810
rect 127906 299730 138822 299810
rect 138994 299730 149910 299810
rect 150082 299730 160998 299810
rect 161170 299730 172086 299810
rect 172258 299730 183174 299810
rect 183346 299730 194262 299810
rect 194434 299730 205350 299810
rect 205522 299730 216438 299810
rect 216610 299730 227526 299810
rect 227698 299730 238614 299810
rect 238786 299730 249702 299810
rect 249874 299730 260790 299810
rect 260962 299730 271878 299810
rect 272050 299730 282966 299810
rect 283138 299730 294054 299810
rect 294226 299730 299250 299810
rect 1246 270 299250 299730
rect 1246 9 6606 270
rect 6778 9 7558 270
rect 7730 9 8510 270
rect 8682 9 9462 270
rect 9634 9 10414 270
rect 10586 9 11366 270
rect 11538 9 12318 270
rect 12490 9 13270 270
rect 13442 9 14222 270
rect 14394 9 15174 270
rect 15346 9 16126 270
rect 16298 9 17078 270
rect 17250 9 18030 270
rect 18202 9 18982 270
rect 19154 9 19934 270
rect 20106 9 20886 270
rect 21058 9 21838 270
rect 22010 9 22790 270
rect 22962 9 23742 270
rect 23914 9 24694 270
rect 24866 9 25646 270
rect 25818 9 26598 270
rect 26770 9 27550 270
rect 27722 9 28502 270
rect 28674 9 29454 270
rect 29626 9 30406 270
rect 30578 9 31358 270
rect 31530 9 32310 270
rect 32482 9 33262 270
rect 33434 9 34214 270
rect 34386 9 35166 270
rect 35338 9 36118 270
rect 36290 9 37070 270
rect 37242 9 38022 270
rect 38194 9 38974 270
rect 39146 9 39926 270
rect 40098 9 40878 270
rect 41050 9 41830 270
rect 42002 9 42782 270
rect 42954 9 43734 270
rect 43906 9 44686 270
rect 44858 9 45638 270
rect 45810 9 46590 270
rect 46762 9 47542 270
rect 47714 9 48494 270
rect 48666 9 49446 270
rect 49618 9 50398 270
rect 50570 9 51350 270
rect 51522 9 52302 270
rect 52474 9 53254 270
rect 53426 9 54206 270
rect 54378 9 55158 270
rect 55330 9 56110 270
rect 56282 9 57062 270
rect 57234 9 58014 270
rect 58186 9 58966 270
rect 59138 9 59918 270
rect 60090 9 60870 270
rect 61042 9 61822 270
rect 61994 9 62774 270
rect 62946 9 63726 270
rect 63898 9 64678 270
rect 64850 9 65630 270
rect 65802 9 66582 270
rect 66754 9 67534 270
rect 67706 9 68486 270
rect 68658 9 69438 270
rect 69610 9 70390 270
rect 70562 9 71342 270
rect 71514 9 72294 270
rect 72466 9 73246 270
rect 73418 9 74198 270
rect 74370 9 75150 270
rect 75322 9 76102 270
rect 76274 9 77054 270
rect 77226 9 78006 270
rect 78178 9 78958 270
rect 79130 9 79910 270
rect 80082 9 80862 270
rect 81034 9 81814 270
rect 81986 9 82766 270
rect 82938 9 83718 270
rect 83890 9 84670 270
rect 84842 9 85622 270
rect 85794 9 86574 270
rect 86746 9 87526 270
rect 87698 9 88478 270
rect 88650 9 89430 270
rect 89602 9 90382 270
rect 90554 9 91334 270
rect 91506 9 92286 270
rect 92458 9 93238 270
rect 93410 9 94190 270
rect 94362 9 95142 270
rect 95314 9 96094 270
rect 96266 9 97046 270
rect 97218 9 97998 270
rect 98170 9 98950 270
rect 99122 9 99902 270
rect 100074 9 100854 270
rect 101026 9 101806 270
rect 101978 9 102758 270
rect 102930 9 103710 270
rect 103882 9 104662 270
rect 104834 9 105614 270
rect 105786 9 106566 270
rect 106738 9 107518 270
rect 107690 9 108470 270
rect 108642 9 109422 270
rect 109594 9 110374 270
rect 110546 9 111326 270
rect 111498 9 112278 270
rect 112450 9 113230 270
rect 113402 9 114182 270
rect 114354 9 115134 270
rect 115306 9 116086 270
rect 116258 9 117038 270
rect 117210 9 117990 270
rect 118162 9 118942 270
rect 119114 9 119894 270
rect 120066 9 120846 270
rect 121018 9 121798 270
rect 121970 9 122750 270
rect 122922 9 123702 270
rect 123874 9 124654 270
rect 124826 9 125606 270
rect 125778 9 126558 270
rect 126730 9 127510 270
rect 127682 9 128462 270
rect 128634 9 129414 270
rect 129586 9 130366 270
rect 130538 9 131318 270
rect 131490 9 132270 270
rect 132442 9 133222 270
rect 133394 9 134174 270
rect 134346 9 135126 270
rect 135298 9 136078 270
rect 136250 9 137030 270
rect 137202 9 137982 270
rect 138154 9 138934 270
rect 139106 9 139886 270
rect 140058 9 140838 270
rect 141010 9 141790 270
rect 141962 9 142742 270
rect 142914 9 143694 270
rect 143866 9 144646 270
rect 144818 9 145598 270
rect 145770 9 146550 270
rect 146722 9 147502 270
rect 147674 9 148454 270
rect 148626 9 149406 270
rect 149578 9 150358 270
rect 150530 9 151310 270
rect 151482 9 152262 270
rect 152434 9 153214 270
rect 153386 9 154166 270
rect 154338 9 155118 270
rect 155290 9 156070 270
rect 156242 9 157022 270
rect 157194 9 157974 270
rect 158146 9 158926 270
rect 159098 9 159878 270
rect 160050 9 160830 270
rect 161002 9 161782 270
rect 161954 9 162734 270
rect 162906 9 163686 270
rect 163858 9 164638 270
rect 164810 9 165590 270
rect 165762 9 166542 270
rect 166714 9 167494 270
rect 167666 9 168446 270
rect 168618 9 169398 270
rect 169570 9 170350 270
rect 170522 9 171302 270
rect 171474 9 172254 270
rect 172426 9 173206 270
rect 173378 9 174158 270
rect 174330 9 175110 270
rect 175282 9 176062 270
rect 176234 9 177014 270
rect 177186 9 177966 270
rect 178138 9 178918 270
rect 179090 9 179870 270
rect 180042 9 180822 270
rect 180994 9 181774 270
rect 181946 9 182726 270
rect 182898 9 183678 270
rect 183850 9 184630 270
rect 184802 9 185582 270
rect 185754 9 186534 270
rect 186706 9 187486 270
rect 187658 9 188438 270
rect 188610 9 189390 270
rect 189562 9 190342 270
rect 190514 9 191294 270
rect 191466 9 192246 270
rect 192418 9 193198 270
rect 193370 9 194150 270
rect 194322 9 195102 270
rect 195274 9 196054 270
rect 196226 9 197006 270
rect 197178 9 197958 270
rect 198130 9 198910 270
rect 199082 9 199862 270
rect 200034 9 200814 270
rect 200986 9 201766 270
rect 201938 9 202718 270
rect 202890 9 203670 270
rect 203842 9 204622 270
rect 204794 9 205574 270
rect 205746 9 206526 270
rect 206698 9 207478 270
rect 207650 9 208430 270
rect 208602 9 209382 270
rect 209554 9 210334 270
rect 210506 9 211286 270
rect 211458 9 212238 270
rect 212410 9 213190 270
rect 213362 9 214142 270
rect 214314 9 215094 270
rect 215266 9 216046 270
rect 216218 9 216998 270
rect 217170 9 217950 270
rect 218122 9 218902 270
rect 219074 9 219854 270
rect 220026 9 220806 270
rect 220978 9 221758 270
rect 221930 9 222710 270
rect 222882 9 223662 270
rect 223834 9 224614 270
rect 224786 9 225566 270
rect 225738 9 226518 270
rect 226690 9 227470 270
rect 227642 9 228422 270
rect 228594 9 229374 270
rect 229546 9 230326 270
rect 230498 9 231278 270
rect 231450 9 232230 270
rect 232402 9 233182 270
rect 233354 9 234134 270
rect 234306 9 235086 270
rect 235258 9 236038 270
rect 236210 9 236990 270
rect 237162 9 237942 270
rect 238114 9 238894 270
rect 239066 9 239846 270
rect 240018 9 240798 270
rect 240970 9 241750 270
rect 241922 9 242702 270
rect 242874 9 243654 270
rect 243826 9 244606 270
rect 244778 9 245558 270
rect 245730 9 246510 270
rect 246682 9 247462 270
rect 247634 9 248414 270
rect 248586 9 249366 270
rect 249538 9 250318 270
rect 250490 9 251270 270
rect 251442 9 252222 270
rect 252394 9 253174 270
rect 253346 9 254126 270
rect 254298 9 255078 270
rect 255250 9 256030 270
rect 256202 9 256982 270
rect 257154 9 257934 270
rect 258106 9 258886 270
rect 259058 9 259838 270
rect 260010 9 260790 270
rect 260962 9 261742 270
rect 261914 9 262694 270
rect 262866 9 263646 270
rect 263818 9 264598 270
rect 264770 9 265550 270
rect 265722 9 266502 270
rect 266674 9 267454 270
rect 267626 9 268406 270
rect 268578 9 269358 270
rect 269530 9 270310 270
rect 270482 9 271262 270
rect 271434 9 272214 270
rect 272386 9 273166 270
rect 273338 9 274118 270
rect 274290 9 275070 270
rect 275242 9 276022 270
rect 276194 9 276974 270
rect 277146 9 277926 270
rect 278098 9 278878 270
rect 279050 9 279830 270
rect 280002 9 280782 270
rect 280954 9 281734 270
rect 281906 9 282686 270
rect 282858 9 283638 270
rect 283810 9 284590 270
rect 284762 9 285542 270
rect 285714 9 286494 270
rect 286666 9 287446 270
rect 287618 9 288398 270
rect 288570 9 289350 270
rect 289522 9 290302 270
rect 290474 9 291254 270
rect 291426 9 292206 270
rect 292378 9 293158 270
rect 293330 9 299250 270
<< metal3 >>
rect 299760 296548 300480 296660
rect -480 295708 240 295820
rect 299760 289884 300480 289996
rect -480 288596 240 288708
rect 299760 283220 300480 283332
rect -480 281484 240 281596
rect 299760 276556 300480 276668
rect -480 274372 240 274484
rect 299760 269892 300480 270004
rect -480 267260 240 267372
rect 299760 263228 300480 263340
rect -480 260148 240 260260
rect 299760 256564 300480 256676
rect -480 253036 240 253148
rect 299760 249900 300480 250012
rect -480 245924 240 246036
rect 299760 243236 300480 243348
rect -480 238812 240 238924
rect 299760 236572 300480 236684
rect -480 231700 240 231812
rect 299760 229908 300480 230020
rect -480 224588 240 224700
rect 299760 223244 300480 223356
rect -480 217476 240 217588
rect 299760 216580 300480 216692
rect -480 210364 240 210476
rect 299760 209916 300480 210028
rect -480 203252 240 203364
rect 299760 203252 300480 203364
rect 299760 196588 300480 196700
rect -480 196140 240 196252
rect 299760 189924 300480 190036
rect -480 189028 240 189140
rect 299760 183260 300480 183372
rect -480 181916 240 182028
rect 299760 176596 300480 176708
rect -480 174804 240 174916
rect 299760 169932 300480 170044
rect -480 167692 240 167804
rect 299760 163268 300480 163380
rect -480 160580 240 160692
rect 299760 156604 300480 156716
rect -480 153468 240 153580
rect 299760 149940 300480 150052
rect -480 146356 240 146468
rect 299760 143276 300480 143388
rect -480 139244 240 139356
rect 299760 136612 300480 136724
rect -480 132132 240 132244
rect 299760 129948 300480 130060
rect -480 125020 240 125132
rect 299760 123284 300480 123396
rect -480 117908 240 118020
rect 299760 116620 300480 116732
rect -480 110796 240 110908
rect 299760 109956 300480 110068
rect -480 103684 240 103796
rect 299760 103292 300480 103404
rect -480 96572 240 96684
rect 299760 96628 300480 96740
rect 299760 89964 300480 90076
rect -480 89460 240 89572
rect 299760 83300 300480 83412
rect -480 82348 240 82460
rect 299760 76636 300480 76748
rect -480 75236 240 75348
rect 299760 69972 300480 70084
rect -480 68124 240 68236
rect 299760 63308 300480 63420
rect -480 61012 240 61124
rect 299760 56644 300480 56756
rect -480 53900 240 54012
rect 299760 49980 300480 50092
rect -480 46788 240 46900
rect 299760 43316 300480 43428
rect -480 39676 240 39788
rect 299760 36652 300480 36764
rect -480 32564 240 32676
rect 299760 29988 300480 30100
rect -480 25452 240 25564
rect 299760 23324 300480 23436
rect -480 18340 240 18452
rect 299760 16660 300480 16772
rect -480 11228 240 11340
rect 299760 9996 300480 10108
rect -480 4116 240 4228
rect 299760 3332 300480 3444
<< obsm3 >>
rect 182 296690 299810 297906
rect 182 296518 299730 296690
rect 182 295850 299810 296518
rect 270 295678 299810 295850
rect 182 290026 299810 295678
rect 182 289854 299730 290026
rect 182 288738 299810 289854
rect 270 288566 299810 288738
rect 182 283362 299810 288566
rect 182 283190 299730 283362
rect 182 281626 299810 283190
rect 270 281454 299810 281626
rect 182 276698 299810 281454
rect 182 276526 299730 276698
rect 182 274514 299810 276526
rect 270 274342 299810 274514
rect 182 270034 299810 274342
rect 182 269862 299730 270034
rect 182 267402 299810 269862
rect 270 267230 299810 267402
rect 182 263370 299810 267230
rect 182 263198 299730 263370
rect 182 260290 299810 263198
rect 270 260118 299810 260290
rect 182 256706 299810 260118
rect 182 256534 299730 256706
rect 182 253178 299810 256534
rect 270 253006 299810 253178
rect 182 250042 299810 253006
rect 182 249870 299730 250042
rect 182 246066 299810 249870
rect 270 245894 299810 246066
rect 182 243378 299810 245894
rect 182 243206 299730 243378
rect 182 238954 299810 243206
rect 270 238782 299810 238954
rect 182 236714 299810 238782
rect 182 236542 299730 236714
rect 182 231842 299810 236542
rect 270 231670 299810 231842
rect 182 230050 299810 231670
rect 182 229878 299730 230050
rect 182 224730 299810 229878
rect 270 224558 299810 224730
rect 182 223386 299810 224558
rect 182 223214 299730 223386
rect 182 217618 299810 223214
rect 270 217446 299810 217618
rect 182 216722 299810 217446
rect 182 216550 299730 216722
rect 182 210506 299810 216550
rect 270 210334 299810 210506
rect 182 210058 299810 210334
rect 182 209886 299730 210058
rect 182 203394 299810 209886
rect 270 203222 299730 203394
rect 182 196730 299810 203222
rect 182 196558 299730 196730
rect 182 196282 299810 196558
rect 270 196110 299810 196282
rect 182 190066 299810 196110
rect 182 189894 299730 190066
rect 182 189170 299810 189894
rect 270 188998 299810 189170
rect 182 183402 299810 188998
rect 182 183230 299730 183402
rect 182 182058 299810 183230
rect 270 181886 299810 182058
rect 182 176738 299810 181886
rect 182 176566 299730 176738
rect 182 174946 299810 176566
rect 270 174774 299810 174946
rect 182 170074 299810 174774
rect 182 169902 299730 170074
rect 182 167834 299810 169902
rect 270 167662 299810 167834
rect 182 163410 299810 167662
rect 182 163238 299730 163410
rect 182 160722 299810 163238
rect 270 160550 299810 160722
rect 182 156746 299810 160550
rect 182 156574 299730 156746
rect 182 153610 299810 156574
rect 270 153438 299810 153610
rect 182 150082 299810 153438
rect 182 149910 299730 150082
rect 182 146498 299810 149910
rect 270 146326 299810 146498
rect 182 143418 299810 146326
rect 182 143246 299730 143418
rect 182 139386 299810 143246
rect 270 139214 299810 139386
rect 182 136754 299810 139214
rect 182 136582 299730 136754
rect 182 132274 299810 136582
rect 270 132102 299810 132274
rect 182 130090 299810 132102
rect 182 129918 299730 130090
rect 182 125162 299810 129918
rect 270 124990 299810 125162
rect 182 123426 299810 124990
rect 182 123254 299730 123426
rect 182 118050 299810 123254
rect 270 117878 299810 118050
rect 182 116762 299810 117878
rect 182 116590 299730 116762
rect 182 110938 299810 116590
rect 270 110766 299810 110938
rect 182 110098 299810 110766
rect 182 109926 299730 110098
rect 182 103826 299810 109926
rect 270 103654 299810 103826
rect 182 103434 299810 103654
rect 182 103262 299730 103434
rect 182 96770 299810 103262
rect 182 96714 299730 96770
rect 270 96598 299730 96714
rect 270 96542 299810 96598
rect 182 90106 299810 96542
rect 182 89934 299730 90106
rect 182 89602 299810 89934
rect 270 89430 299810 89602
rect 182 83442 299810 89430
rect 182 83270 299730 83442
rect 182 82490 299810 83270
rect 270 82318 299810 82490
rect 182 76778 299810 82318
rect 182 76606 299730 76778
rect 182 75378 299810 76606
rect 270 75206 299810 75378
rect 182 70114 299810 75206
rect 182 69942 299730 70114
rect 182 68266 299810 69942
rect 270 68094 299810 68266
rect 182 63450 299810 68094
rect 182 63278 299730 63450
rect 182 61154 299810 63278
rect 270 60982 299810 61154
rect 182 56786 299810 60982
rect 182 56614 299730 56786
rect 182 54042 299810 56614
rect 270 53870 299810 54042
rect 182 50122 299810 53870
rect 182 49950 299730 50122
rect 182 46930 299810 49950
rect 270 46758 299810 46930
rect 182 43458 299810 46758
rect 182 43286 299730 43458
rect 182 39818 299810 43286
rect 270 39646 299810 39818
rect 182 36794 299810 39646
rect 182 36622 299730 36794
rect 182 32706 299810 36622
rect 270 32534 299810 32706
rect 182 30130 299810 32534
rect 182 29958 299730 30130
rect 182 25594 299810 29958
rect 270 25422 299810 25594
rect 182 23466 299810 25422
rect 182 23294 299730 23466
rect 182 18482 299810 23294
rect 270 18310 299810 18482
rect 182 16802 299810 18310
rect 182 16630 299730 16802
rect 182 11370 299810 16630
rect 270 11198 299810 11370
rect 182 10138 299810 11198
rect 182 9966 299730 10138
rect 182 4258 299810 9966
rect 270 4086 299810 4258
rect 182 3474 299810 4086
rect 182 3302 299730 3474
rect 182 14 299810 3302
<< metal4 >>
rect -6 162 304 299718
rect 474 642 784 299238
rect 2529 162 2839 299718
rect 4389 162 4699 299718
rect 11529 162 11839 299718
rect 13389 162 13699 299718
rect 20529 162 20839 299718
rect 22389 162 22699 299718
rect 29529 162 29839 299718
rect 31389 162 31699 299718
rect 38529 162 38839 299718
rect 40389 162 40699 299718
rect 47529 162 47839 299718
rect 49389 162 49699 299718
rect 56529 162 56839 299718
rect 58389 162 58699 299718
rect 65529 162 65839 299718
rect 67389 162 67699 299718
rect 74529 162 74839 299718
rect 76389 162 76699 299718
rect 83529 162 83839 299718
rect 85389 162 85699 299718
rect 92529 162 92839 299718
rect 94389 162 94699 299718
rect 101529 162 101839 299718
rect 103389 134458 103699 299718
rect 103389 162 103699 55510
rect 110529 162 110839 299718
rect 112389 162 112699 299718
rect 119529 162 119839 299718
rect 121389 162 121699 299718
rect 128529 162 128839 299718
rect 130389 162 130699 299718
rect 137529 162 137839 299718
rect 139389 162 139699 299718
rect 146529 162 146839 299718
rect 148389 162 148699 299718
rect 155529 162 155839 299718
rect 157389 162 157699 299718
rect 164529 162 164839 299718
rect 166389 162 166699 299718
rect 173529 162 173839 299718
rect 175389 162 175699 299718
rect 182529 162 182839 299718
rect 184389 162 184699 299718
rect 191529 162 191839 299718
rect 193389 162 193699 299718
rect 200529 162 200839 299718
rect 202389 162 202699 299718
rect 209529 162 209839 299718
rect 211389 162 211699 299718
rect 218529 162 218839 299718
rect 220389 162 220699 299718
rect 227529 162 227839 299718
rect 229389 162 229699 299718
rect 236529 162 236839 299718
rect 238389 162 238699 299718
rect 245529 162 245839 299718
rect 247389 162 247699 299718
rect 254529 162 254839 299718
rect 256389 162 256699 299718
rect 263529 162 263839 299718
rect 265389 162 265699 299718
rect 272529 162 272839 299718
rect 274389 162 274699 299718
rect 281529 162 281839 299718
rect 283389 162 283699 299718
rect 290529 162 290839 299718
rect 292389 162 292699 299718
rect 299208 642 299518 299238
rect 299688 162 299998 299718
<< obsm4 >>
rect 39886 2025 40359 297855
rect 40729 2025 47499 297855
rect 47869 2025 49359 297855
rect 49729 2025 56499 297855
rect 56869 2025 58359 297855
rect 58729 2025 65499 297855
rect 65869 2025 67359 297855
rect 67729 2025 74499 297855
rect 74869 2025 76359 297855
rect 76729 2025 83499 297855
rect 83869 2025 85359 297855
rect 85729 2025 92499 297855
rect 92869 2025 94359 297855
rect 94729 2025 101499 297855
rect 101869 134428 103359 297855
rect 103729 134428 110499 297855
rect 101869 55540 110499 134428
rect 101869 2025 103359 55540
rect 103729 2025 110499 55540
rect 110869 2025 112359 297855
rect 112729 2025 119499 297855
rect 119869 2025 121359 297855
rect 121729 2025 128499 297855
rect 128869 2025 130359 297855
rect 130729 2025 137499 297855
rect 137869 2025 139359 297855
rect 139729 2025 146499 297855
rect 146869 2025 148359 297855
rect 148729 2025 150122 297855
<< metal5 >>
rect -6 299408 299998 299718
rect 474 298928 299518 299238
rect -6 293697 299998 294007
rect -6 290697 299998 291007
rect -6 284697 299998 285007
rect -6 281697 299998 282007
rect -6 275697 299998 276007
rect -6 272697 299998 273007
rect -6 266697 299998 267007
rect -6 263697 299998 264007
rect -6 257697 299998 258007
rect -6 254697 299998 255007
rect -6 248697 299998 249007
rect -6 245697 299998 246007
rect -6 239697 299998 240007
rect -6 236697 299998 237007
rect -6 230697 299998 231007
rect -6 227697 299998 228007
rect -6 221697 299998 222007
rect -6 218697 299998 219007
rect -6 212697 299998 213007
rect -6 209697 299998 210007
rect -6 203697 299998 204007
rect -6 200697 299998 201007
rect -6 194697 299998 195007
rect -6 191697 299998 192007
rect -6 185697 299998 186007
rect -6 182697 299998 183007
rect -6 176697 299998 177007
rect -6 173697 299998 174007
rect -6 167697 299998 168007
rect -6 164697 299998 165007
rect -6 158697 299998 159007
rect -6 155697 299998 156007
rect -6 149697 299998 150007
rect -6 146697 299998 147007
rect -6 140697 299998 141007
rect -6 137697 299998 138007
rect -6 131697 299998 132007
rect -6 128697 299998 129007
rect -6 122697 299998 123007
rect -6 119697 299998 120007
rect -6 113697 299998 114007
rect -6 110697 299998 111007
rect -6 104697 299998 105007
rect -6 101697 299998 102007
rect -6 95697 299998 96007
rect -6 92697 299998 93007
rect -6 86697 299998 87007
rect -6 83697 299998 84007
rect -6 77697 299998 78007
rect -6 74697 299998 75007
rect -6 68697 299998 69007
rect -6 65697 299998 66007
rect -6 59697 299998 60007
rect -6 56697 299998 57007
rect -6 50697 299998 51007
rect -6 47697 299998 48007
rect -6 41697 299998 42007
rect -6 38697 299998 39007
rect -6 32697 299998 33007
rect -6 29697 299998 30007
rect -6 23697 299998 24007
rect -6 20697 299998 21007
rect -6 14697 299998 15007
rect -6 11697 299998 12007
rect -6 5697 299998 6007
rect -6 2697 299998 3007
rect 474 642 299518 952
rect -6 162 299998 472
<< labels >>
rlabel metal3 s 299760 3332 300480 3444 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 299760 203252 300480 203364 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 299760 223244 300480 223356 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 299760 243236 300480 243348 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 299760 263228 300480 263340 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 299760 283220 300480 283332 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 294084 299760 294196 300480 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 260820 299760 260932 300480 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 227556 299760 227668 300480 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 194292 299760 194404 300480 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 161028 299760 161140 300480 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 299760 23324 300480 23436 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 127764 299760 127876 300480 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 94500 299760 94612 300480 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 61236 299760 61348 300480 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 27972 299760 28084 300480 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s -480 295708 240 295820 4 io_in[24]
port 17 nsew signal input
rlabel metal3 s -480 274372 240 274484 4 io_in[25]
port 18 nsew signal input
rlabel metal3 s -480 253036 240 253148 4 io_in[26]
port 19 nsew signal input
rlabel metal3 s -480 231700 240 231812 4 io_in[27]
port 20 nsew signal input
rlabel metal3 s -480 210364 240 210476 4 io_in[28]
port 21 nsew signal input
rlabel metal3 s -480 189028 240 189140 4 io_in[29]
port 22 nsew signal input
rlabel metal3 s 299760 43316 300480 43428 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s -480 167692 240 167804 4 io_in[30]
port 24 nsew signal input
rlabel metal3 s -480 146356 240 146468 4 io_in[31]
port 25 nsew signal input
rlabel metal3 s -480 125020 240 125132 4 io_in[32]
port 26 nsew signal input
rlabel metal3 s -480 103684 240 103796 4 io_in[33]
port 27 nsew signal input
rlabel metal3 s -480 82348 240 82460 4 io_in[34]
port 28 nsew signal input
rlabel metal3 s -480 61012 240 61124 4 io_in[35]
port 29 nsew signal input
rlabel metal3 s -480 39676 240 39788 4 io_in[36]
port 30 nsew signal input
rlabel metal3 s -480 18340 240 18452 4 io_in[37]
port 31 nsew signal input
rlabel metal3 s 299760 63308 300480 63420 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 299760 83300 300480 83412 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 299760 103292 300480 103404 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 299760 123284 300480 123396 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 299760 143276 300480 143388 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 299760 163268 300480 163380 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 299760 183260 300480 183372 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 299760 16660 300480 16772 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 299760 216580 300480 216692 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 299760 236572 300480 236684 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 299760 256564 300480 256676 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 299760 276556 300480 276668 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 299760 296548 300480 296660 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 271908 299760 272020 300480 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 238644 299760 238756 300480 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 205380 299760 205492 300480 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 172116 299760 172228 300480 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 138852 299760 138964 300480 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 299760 36652 300480 36764 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 105588 299760 105700 300480 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 72324 299760 72436 300480 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 39060 299760 39172 300480 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 5796 299760 5908 300480 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s -480 281484 240 281596 4 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s -480 260148 240 260260 4 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s -480 238812 240 238924 4 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s -480 217476 240 217588 4 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s -480 196140 240 196252 4 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s -480 174804 240 174916 4 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 299760 56644 300480 56756 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s -480 153468 240 153580 4 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s -480 132132 240 132244 4 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s -480 110796 240 110908 4 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s -480 89460 240 89572 4 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s -480 68124 240 68236 4 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s -480 46788 240 46900 4 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s -480 25452 240 25564 4 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s -480 4116 240 4228 4 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 299760 76636 300480 76748 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 299760 96628 300480 96740 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 299760 116620 300480 116732 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 299760 136612 300480 136724 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 299760 156604 300480 156716 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 299760 176596 300480 176708 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 299760 196588 300480 196700 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 299760 9996 300480 10108 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 299760 209916 300480 210028 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 299760 229908 300480 230020 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 299760 249900 300480 250012 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 299760 269892 300480 270004 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 299760 289884 300480 289996 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 282996 299760 283108 300480 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 249732 299760 249844 300480 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 216468 299760 216580 300480 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 183204 299760 183316 300480 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 149940 299760 150052 300480 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 299760 29988 300480 30100 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 116676 299760 116788 300480 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 83412 299760 83524 300480 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 50148 299760 50260 300480 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 16884 299760 16996 300480 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s -480 288596 240 288708 4 io_out[24]
port 93 nsew signal output
rlabel metal3 s -480 267260 240 267372 4 io_out[25]
port 94 nsew signal output
rlabel metal3 s -480 245924 240 246036 4 io_out[26]
port 95 nsew signal output
rlabel metal3 s -480 224588 240 224700 4 io_out[27]
port 96 nsew signal output
rlabel metal3 s -480 203252 240 203364 4 io_out[28]
port 97 nsew signal output
rlabel metal3 s -480 181916 240 182028 4 io_out[29]
port 98 nsew signal output
rlabel metal3 s 299760 49980 300480 50092 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s -480 160580 240 160692 4 io_out[30]
port 100 nsew signal output
rlabel metal3 s -480 139244 240 139356 4 io_out[31]
port 101 nsew signal output
rlabel metal3 s -480 117908 240 118020 4 io_out[32]
port 102 nsew signal output
rlabel metal3 s -480 96572 240 96684 4 io_out[33]
port 103 nsew signal output
rlabel metal3 s -480 75236 240 75348 4 io_out[34]
port 104 nsew signal output
rlabel metal3 s -480 53900 240 54012 4 io_out[35]
port 105 nsew signal output
rlabel metal3 s -480 32564 240 32676 4 io_out[36]
port 106 nsew signal output
rlabel metal3 s -480 11228 240 11340 4 io_out[37]
port 107 nsew signal output
rlabel metal3 s 299760 69972 300480 70084 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 299760 89964 300480 90076 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 299760 109956 300480 110068 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 299760 129948 300480 130060 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 299760 149940 300480 150052 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 299760 169932 300480 170044 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 299760 189924 300480 190036 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 107548 -480 107660 240 8 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 136108 -480 136220 240 8 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 138964 -480 139076 240 8 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 141820 -480 141932 240 8 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 144676 -480 144788 240 8 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 147532 -480 147644 240 8 la_data_in[14]
port 120 nsew signal input
rlabel metal2 s 150388 -480 150500 240 8 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 153244 -480 153356 240 8 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 156100 -480 156212 240 8 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 158956 -480 159068 240 8 la_data_in[18]
port 124 nsew signal input
rlabel metal2 s 161812 -480 161924 240 8 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 110404 -480 110516 240 8 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 164668 -480 164780 240 8 la_data_in[20]
port 127 nsew signal input
rlabel metal2 s 167524 -480 167636 240 8 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 170380 -480 170492 240 8 la_data_in[22]
port 129 nsew signal input
rlabel metal2 s 173236 -480 173348 240 8 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 176092 -480 176204 240 8 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 178948 -480 179060 240 8 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 181804 -480 181916 240 8 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 184660 -480 184772 240 8 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 187516 -480 187628 240 8 la_data_in[28]
port 135 nsew signal input
rlabel metal2 s 190372 -480 190484 240 8 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 113260 -480 113372 240 8 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 193228 -480 193340 240 8 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 196084 -480 196196 240 8 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 198940 -480 199052 240 8 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 201796 -480 201908 240 8 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 204652 -480 204764 240 8 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 207508 -480 207620 240 8 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 210364 -480 210476 240 8 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 213220 -480 213332 240 8 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 216076 -480 216188 240 8 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 218932 -480 219044 240 8 la_data_in[39]
port 147 nsew signal input
rlabel metal2 s 116116 -480 116228 240 8 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 221788 -480 221900 240 8 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 224644 -480 224756 240 8 la_data_in[41]
port 150 nsew signal input
rlabel metal2 s 227500 -480 227612 240 8 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 230356 -480 230468 240 8 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 233212 -480 233324 240 8 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 236068 -480 236180 240 8 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 238924 -480 239036 240 8 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 241780 -480 241892 240 8 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 244636 -480 244748 240 8 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 247492 -480 247604 240 8 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 118972 -480 119084 240 8 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 250348 -480 250460 240 8 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 253204 -480 253316 240 8 la_data_in[51]
port 161 nsew signal input
rlabel metal2 s 256060 -480 256172 240 8 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 258916 -480 259028 240 8 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 261772 -480 261884 240 8 la_data_in[54]
port 164 nsew signal input
rlabel metal2 s 264628 -480 264740 240 8 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 267484 -480 267596 240 8 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 270340 -480 270452 240 8 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 273196 -480 273308 240 8 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 276052 -480 276164 240 8 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 121828 -480 121940 240 8 la_data_in[5]
port 170 nsew signal input
rlabel metal2 s 278908 -480 279020 240 8 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 281764 -480 281876 240 8 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 284620 -480 284732 240 8 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 287476 -480 287588 240 8 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 124684 -480 124796 240 8 la_data_in[6]
port 175 nsew signal input
rlabel metal2 s 127540 -480 127652 240 8 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 130396 -480 130508 240 8 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 133252 -480 133364 240 8 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 108500 -480 108612 240 8 la_data_out[0]
port 179 nsew signal output
rlabel metal2 s 137060 -480 137172 240 8 la_data_out[10]
port 180 nsew signal output
rlabel metal2 s 139916 -480 140028 240 8 la_data_out[11]
port 181 nsew signal output
rlabel metal2 s 142772 -480 142884 240 8 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 145628 -480 145740 240 8 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 148484 -480 148596 240 8 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 151340 -480 151452 240 8 la_data_out[15]
port 185 nsew signal output
rlabel metal2 s 154196 -480 154308 240 8 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 157052 -480 157164 240 8 la_data_out[17]
port 187 nsew signal output
rlabel metal2 s 159908 -480 160020 240 8 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 162764 -480 162876 240 8 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 111356 -480 111468 240 8 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 165620 -480 165732 240 8 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 168476 -480 168588 240 8 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 171332 -480 171444 240 8 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 174188 -480 174300 240 8 la_data_out[23]
port 194 nsew signal output
rlabel metal2 s 177044 -480 177156 240 8 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 179900 -480 180012 240 8 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 182756 -480 182868 240 8 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 185612 -480 185724 240 8 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 188468 -480 188580 240 8 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 191324 -480 191436 240 8 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 114212 -480 114324 240 8 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 194180 -480 194292 240 8 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 197036 -480 197148 240 8 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 199892 -480 200004 240 8 la_data_out[32]
port 204 nsew signal output
rlabel metal2 s 202748 -480 202860 240 8 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 205604 -480 205716 240 8 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 208460 -480 208572 240 8 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 211316 -480 211428 240 8 la_data_out[36]
port 208 nsew signal output
rlabel metal2 s 214172 -480 214284 240 8 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 217028 -480 217140 240 8 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 219884 -480 219996 240 8 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 117068 -480 117180 240 8 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 222740 -480 222852 240 8 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 225596 -480 225708 240 8 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 228452 -480 228564 240 8 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 231308 -480 231420 240 8 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 234164 -480 234276 240 8 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 237020 -480 237132 240 8 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 239876 -480 239988 240 8 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 242732 -480 242844 240 8 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 245588 -480 245700 240 8 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 248444 -480 248556 240 8 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 119924 -480 120036 240 8 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 251300 -480 251412 240 8 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 254156 -480 254268 240 8 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 257012 -480 257124 240 8 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 259868 -480 259980 240 8 la_data_out[53]
port 227 nsew signal output
rlabel metal2 s 262724 -480 262836 240 8 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 265580 -480 265692 240 8 la_data_out[55]
port 229 nsew signal output
rlabel metal2 s 268436 -480 268548 240 8 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 271292 -480 271404 240 8 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 274148 -480 274260 240 8 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 277004 -480 277116 240 8 la_data_out[59]
port 233 nsew signal output
rlabel metal2 s 122780 -480 122892 240 8 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 279860 -480 279972 240 8 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 282716 -480 282828 240 8 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 285572 -480 285684 240 8 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 288428 -480 288540 240 8 la_data_out[63]
port 238 nsew signal output
rlabel metal2 s 125636 -480 125748 240 8 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 128492 -480 128604 240 8 la_data_out[7]
port 240 nsew signal output
rlabel metal2 s 131348 -480 131460 240 8 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 134204 -480 134316 240 8 la_data_out[9]
port 242 nsew signal output
rlabel metal2 s 109452 -480 109564 240 8 la_oenb[0]
port 243 nsew signal input
rlabel metal2 s 138012 -480 138124 240 8 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 140868 -480 140980 240 8 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 143724 -480 143836 240 8 la_oenb[12]
port 246 nsew signal input
rlabel metal2 s 146580 -480 146692 240 8 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 149436 -480 149548 240 8 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 152292 -480 152404 240 8 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 155148 -480 155260 240 8 la_oenb[16]
port 250 nsew signal input
rlabel metal2 s 158004 -480 158116 240 8 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 160860 -480 160972 240 8 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 163716 -480 163828 240 8 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 112308 -480 112420 240 8 la_oenb[1]
port 254 nsew signal input
rlabel metal2 s 166572 -480 166684 240 8 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 169428 -480 169540 240 8 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 172284 -480 172396 240 8 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 175140 -480 175252 240 8 la_oenb[23]
port 258 nsew signal input
rlabel metal2 s 177996 -480 178108 240 8 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 180852 -480 180964 240 8 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 183708 -480 183820 240 8 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 186564 -480 186676 240 8 la_oenb[27]
port 262 nsew signal input
rlabel metal2 s 189420 -480 189532 240 8 la_oenb[28]
port 263 nsew signal input
rlabel metal2 s 192276 -480 192388 240 8 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 115164 -480 115276 240 8 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 195132 -480 195244 240 8 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 197988 -480 198100 240 8 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 200844 -480 200956 240 8 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 203700 -480 203812 240 8 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 206556 -480 206668 240 8 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 209412 -480 209524 240 8 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 212268 -480 212380 240 8 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 215124 -480 215236 240 8 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 217980 -480 218092 240 8 la_oenb[38]
port 274 nsew signal input
rlabel metal2 s 220836 -480 220948 240 8 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 118020 -480 118132 240 8 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 223692 -480 223804 240 8 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 226548 -480 226660 240 8 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 229404 -480 229516 240 8 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 232260 -480 232372 240 8 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 235116 -480 235228 240 8 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 237972 -480 238084 240 8 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 240828 -480 240940 240 8 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 243684 -480 243796 240 8 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 246540 -480 246652 240 8 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 249396 -480 249508 240 8 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 120876 -480 120988 240 8 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 252252 -480 252364 240 8 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 255108 -480 255220 240 8 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 257964 -480 258076 240 8 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 260820 -480 260932 240 8 la_oenb[53]
port 291 nsew signal input
rlabel metal2 s 263676 -480 263788 240 8 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 266532 -480 266644 240 8 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 269388 -480 269500 240 8 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 272244 -480 272356 240 8 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 275100 -480 275212 240 8 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 277956 -480 278068 240 8 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 123732 -480 123844 240 8 la_oenb[5]
port 298 nsew signal input
rlabel metal2 s 280812 -480 280924 240 8 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 283668 -480 283780 240 8 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 286524 -480 286636 240 8 la_oenb[62]
port 301 nsew signal input
rlabel metal2 s 289380 -480 289492 240 8 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 126588 -480 126700 240 8 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 129444 -480 129556 240 8 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 132300 -480 132412 240 8 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 135156 -480 135268 240 8 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 290332 -480 290444 240 8 user_clock2
port 307 nsew signal input
rlabel metal2 s 291284 -480 291396 240 8 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 292236 -480 292348 240 8 user_irq[1]
port 309 nsew signal output
rlabel metal2 s 293188 -480 293300 240 8 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 474 642 784 299238 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 474 642 299518 952 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s 474 298928 299518 299238 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 299208 642 299518 299238 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 2529 162 2839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 11529 162 11839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 20529 162 20839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 29529 162 29839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 38529 162 38839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 47529 162 47839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 56529 162 56839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 65529 162 65839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 74529 162 74839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 83529 162 83839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 92529 162 92839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 101529 162 101839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 110529 162 110839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 119529 162 119839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 128529 162 128839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 137529 162 137839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 146529 162 146839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 155529 162 155839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 164529 162 164839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 173529 162 173839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 182529 162 182839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 191529 162 191839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 200529 162 200839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 209529 162 209839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 218529 162 218839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 227529 162 227839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 236529 162 236839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 245529 162 245839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 254529 162 254839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 263529 162 263839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 272529 162 272839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 281529 162 281839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 290529 162 290839 299718 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 2697 299998 3007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 11697 299998 12007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 20697 299998 21007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 29697 299998 30007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 38697 299998 39007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 47697 299998 48007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 56697 299998 57007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 65697 299998 66007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 74697 299998 75007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 83697 299998 84007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 92697 299998 93007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 101697 299998 102007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 110697 299998 111007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 119697 299998 120007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 128697 299998 129007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 137697 299998 138007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 146697 299998 147007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 155697 299998 156007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 164697 299998 165007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 173697 299998 174007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 182697 299998 183007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 191697 299998 192007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 200697 299998 201007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 209697 299998 210007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 218697 299998 219007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 227697 299998 228007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 236697 299998 237007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 245697 299998 246007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 254697 299998 255007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 263697 299998 264007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 272697 299998 273007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 281697 299998 282007 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -6 290697 299998 291007 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s -6 162 304 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 162 299998 472 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 299408 299998 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 299688 162 299998 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 4389 162 4699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 13389 162 13699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 22389 162 22699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 31389 162 31699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40389 162 40699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 49389 162 49699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 58389 162 58699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 67389 162 67699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 76389 162 76699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 85389 162 85699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 94389 162 94699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 103389 162 103699 55510 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 103389 134458 103699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 112389 162 112699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 121389 162 121699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 130389 162 130699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 139389 162 139699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 148389 162 148699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 157389 162 157699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 166389 162 166699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 175389 162 175699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 184389 162 184699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 193389 162 193699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 202389 162 202699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 211389 162 211699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 220389 162 220699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 229389 162 229699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 238389 162 238699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 247389 162 247699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 256389 162 256699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 265389 162 265699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 274389 162 274699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 283389 162 283699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 292389 162 292699 299718 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 5697 299998 6007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 14697 299998 15007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 23697 299998 24007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 32697 299998 33007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 41697 299998 42007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 50697 299998 51007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 59697 299998 60007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 68697 299998 69007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 77697 299998 78007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 86697 299998 87007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 95697 299998 96007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 104697 299998 105007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 113697 299998 114007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 122697 299998 123007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 131697 299998 132007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 140697 299998 141007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 149697 299998 150007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 158697 299998 159007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 167697 299998 168007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 176697 299998 177007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 185697 299998 186007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 194697 299998 195007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 203697 299998 204007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 212697 299998 213007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 221697 299998 222007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 230697 299998 231007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 239697 299998 240007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 248697 299998 249007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 257697 299998 258007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 266697 299998 267007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 275697 299998 276007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 284697 299998 285007 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -6 293697 299998 294007 6 vss
port 312 nsew ground bidirectional
rlabel metal2 s 6636 -480 6748 240 8 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 7588 -480 7700 240 8 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 8540 -480 8652 240 8 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 12348 -480 12460 240 8 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 44716 -480 44828 240 8 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 47572 -480 47684 240 8 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 50428 -480 50540 240 8 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 53284 -480 53396 240 8 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 56140 -480 56252 240 8 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 58996 -480 59108 240 8 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 61852 -480 61964 240 8 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 64708 -480 64820 240 8 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 67564 -480 67676 240 8 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 70420 -480 70532 240 8 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 16156 -480 16268 240 8 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 73276 -480 73388 240 8 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 76132 -480 76244 240 8 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 78988 -480 79100 240 8 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 81844 -480 81956 240 8 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 84700 -480 84812 240 8 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 87556 -480 87668 240 8 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 90412 -480 90524 240 8 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 93268 -480 93380 240 8 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 96124 -480 96236 240 8 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 98980 -480 99092 240 8 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 19964 -480 20076 240 8 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 101836 -480 101948 240 8 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 104692 -480 104804 240 8 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 23772 -480 23884 240 8 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 27580 -480 27692 240 8 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 30436 -480 30548 240 8 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 33292 -480 33404 240 8 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 36148 -480 36260 240 8 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 39004 -480 39116 240 8 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 41860 -480 41972 240 8 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 9492 -480 9604 240 8 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 13300 -480 13412 240 8 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 45668 -480 45780 240 8 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 48524 -480 48636 240 8 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 51380 -480 51492 240 8 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 54236 -480 54348 240 8 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 57092 -480 57204 240 8 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 59948 -480 60060 240 8 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 62804 -480 62916 240 8 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 65660 -480 65772 240 8 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 68516 -480 68628 240 8 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 71372 -480 71484 240 8 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 17108 -480 17220 240 8 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 74228 -480 74340 240 8 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 77084 -480 77196 240 8 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 79940 -480 80052 240 8 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 82796 -480 82908 240 8 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 85652 -480 85764 240 8 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 88508 -480 88620 240 8 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 91364 -480 91476 240 8 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 94220 -480 94332 240 8 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 97076 -480 97188 240 8 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 99932 -480 100044 240 8 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 20916 -480 21028 240 8 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 102788 -480 102900 240 8 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 105644 -480 105756 240 8 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 24724 -480 24836 240 8 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 28532 -480 28644 240 8 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 31388 -480 31500 240 8 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 34244 -480 34356 240 8 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 37100 -480 37212 240 8 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 39956 -480 40068 240 8 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 42812 -480 42924 240 8 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 14252 -480 14364 240 8 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 46620 -480 46732 240 8 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 49476 -480 49588 240 8 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 52332 -480 52444 240 8 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 55188 -480 55300 240 8 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 58044 -480 58156 240 8 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 60900 -480 61012 240 8 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 63756 -480 63868 240 8 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 66612 -480 66724 240 8 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 69468 -480 69580 240 8 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 72324 -480 72436 240 8 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 18060 -480 18172 240 8 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 75180 -480 75292 240 8 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 78036 -480 78148 240 8 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 80892 -480 81004 240 8 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 83748 -480 83860 240 8 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 86604 -480 86716 240 8 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 89460 -480 89572 240 8 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 92316 -480 92428 240 8 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 95172 -480 95284 240 8 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 98028 -480 98140 240 8 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 100884 -480 100996 240 8 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 21868 -480 21980 240 8 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 103740 -480 103852 240 8 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 106596 -480 106708 240 8 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 25676 -480 25788 240 8 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 29484 -480 29596 240 8 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 32340 -480 32452 240 8 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 35196 -480 35308 240 8 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 38052 -480 38164 240 8 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 40908 -480 41020 240 8 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 43764 -480 43876 240 8 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 15204 -480 15316 240 8 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 19012 -480 19124 240 8 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 22820 -480 22932 240 8 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 26628 -480 26740 240 8 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 10444 -480 10556 240 8 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 11396 -480 11508 240 8 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6329678
string GDS_FILE /home/runner/work/tiny_silicon_1/tiny_silicon_1/openlane/user_project_wrapper/runs/22_12_02_06_06/results/signoff/user_project_wrapper.magic.gds
string GDS_START 3247320
<< end >>

