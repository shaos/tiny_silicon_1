VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 800.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 655.200 4.000 655.760 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 665.280 4.000 665.840 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 325.920 4.000 326.480 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 574.560 4.000 575.120 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 393.120 4.000 393.680 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 336.000 4.000 336.560 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 796.000 652.400 799.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 40.320 1099.000 40.880 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 742.560 1099.000 743.120 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 796.000 790.160 799.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 930.720 1.000 931.280 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 796.000 269.360 799.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 796.000 907.760 799.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 1.000 665.840 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1098.720 796.000 1099.280 799.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 668.640 1099.000 669.200 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 1.000 786.800 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 1.000 128.240 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 792.960 4.000 793.520 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 648.480 4.000 649.040 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 739.200 4.000 739.760 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 591.360 4.000 591.920 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 789.600 1099.000 790.160 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 1.000 622.160 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 399.840 4.000 400.400 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 1.000 803.600 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 97.440 4.000 98.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 796.000 50.960 799.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1001.280 796.000 1001.840 799.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 688.800 1099.000 689.360 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 567.840 1099.000 568.400 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 779.520 1099.000 780.080 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 275.520 1099.000 276.080 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 181.440 4.000 182.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 30.240 1099.000 30.800 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 796.000 927.920 799.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 436.800 4.000 437.360 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 490.560 4.000 491.120 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 514.080 1099.000 514.640 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 460.320 1099.000 460.880 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 796.000 185.360 799.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 1.000 585.200 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 245.280 4.000 245.840 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 1.000 867.440 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 796.000 753.200 799.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 1.000 272.720 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 1.000 91.280 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 796.000 195.440 799.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 796.000 487.760 799.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 796.000 407.120 799.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 796.000 699.440 799.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 1.000 813.680 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 94.080 1099.000 94.640 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1071.840 796.000 1072.400 799.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 272.160 4.000 272.720 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 134.400 4.000 134.960 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 796.000 67.760 799.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 792.960 1.000 793.520 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 796.000 168.560 799.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 332.640 1099.000 333.200 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 211.680 1099.000 212.240 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 893.760 1.000 894.320 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 292.320 4.000 292.880 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 796.000 981.680 799.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 3.360 1099.000 3.920 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 776.160 4.000 776.720 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 705.600 1099.000 706.160 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 796.000 679.280 799.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 231.840 1099.000 232.400 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 712.320 4.000 712.880 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 127.680 4.000 128.240 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 796.000 843.920 799.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 749.280 4.000 749.840 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 796.000 608.720 799.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 473.760 4.000 474.320 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 769.440 1099.000 770.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 796.000 306.320 799.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 796.000 444.080 799.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 1.000 612.080 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1081.920 796.000 1082.480 799.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 796.000 148.400 799.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 702.240 4.000 702.800 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 1.000 383.600 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 641.760 1099.000 642.320 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 1.000 108.080 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 1.000 884.240 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 796.000 360.080 799.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 1.000 64.400 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1041.600 1.000 1042.160 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 628.320 4.000 628.880 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 57.120 1099.000 57.680 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 356.160 4.000 356.720 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 1.000 830.480 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 977.760 1.000 978.320 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 1.000 400.400 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 1.000 319.760 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 796.000 817.040 799.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 1.000 649.040 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 184.800 1099.000 185.360 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 796.000 1018.640 799.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 1.000 336.560 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 796.000 743.120 799.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 346.080 4.000 346.640 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 1.000 628.880 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 1.000 565.040 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 1.000 229.040 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 43.680 4.000 44.240 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 796.000 588.560 799.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 1.000 437.360 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 796.000 551.600 799.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 171.360 4.000 171.920 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 537.600 4.000 538.160 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 1.000 692.720 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 1.000 245.840 4.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 483.840 4.000 484.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 732.480 1099.000 733.040 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 268.800 1099.000 269.360 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 1.000 292.880 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 796.000 534.800 799.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 796.000 30.800 799.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 534.240 1099.000 534.800 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 796.000 242.480 799.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 1.000 1095.920 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 796.000 625.520 799.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 144.480 4.000 145.040 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 796.000 370.160 799.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 47.040 1099.000 47.600 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 719.040 4.000 719.600 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 420.000 4.000 420.560 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 561.120 1099.000 561.680 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 796.000 635.600 799.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 796.000 350.000 799.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 796.000 736.400 799.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 796.000 57.680 799.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 796.000 94.640 799.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 84.000 1099.000 84.560 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 796.000 571.760 799.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 70.560 4.000 71.120 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 796.000 954.800 799.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 383.040 4.000 383.600 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 638.400 4.000 638.960 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 796.000 222.320 799.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 796.000 40.880 799.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 1.000 675.920 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 796.000 131.600 799.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 1.000 427.280 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 796.000 672.560 799.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 369.600 1099.000 370.160 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 1.000 326.480 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 1.000 457.520 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 319.200 4.000 319.760 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1044.960 796.000 1045.520 799.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 1.000 958.160 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 1.000 309.680 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 540.960 1099.000 541.520 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 1.000 591.920 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 796.000 598.640 799.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 796.000 514.640 799.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 796.000 232.400 799.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 796.000 524.720 799.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 446.880 1.000 447.440 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 168.000 1099.000 168.560 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 796.000 890.960 799.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 826.560 796.000 827.120 799.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 255.360 4.000 255.920 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 282.240 4.000 282.800 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 796.000 178.640 799.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 1.000 346.640 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 715.680 1099.000 716.240 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 1.000 161.840 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 477.120 1099.000 477.680 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.880 4.000 27.440 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 1.000 554.960 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 796.000 397.040 799.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 1.000 192.080 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 194.880 1099.000 195.440 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 16.800 4.000 17.360 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1008.000 796.000 1008.560 799.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 796.000 971.600 799.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 359.520 1099.000 360.080 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 33.600 4.000 34.160 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 685.440 4.000 686.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1.000 356.720 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 241.920 1099.000 242.480 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 796.000 14.000 799.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 376.320 1099.000 376.880 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 796.000 615.440 799.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 635.040 1099.000 635.600 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 1.000 501.200 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 295.680 1099.000 296.240 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1085.280 1.000 1085.840 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 796.000 141.680 799.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 440.160 1099.000 440.720 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 1.000 282.800 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 426.720 4.000 427.280 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 1.000 511.280 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 796.000 121.520 799.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 796.000 726.320 799.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 604.800 1099.000 605.360 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 1.000 410.480 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 218.400 4.000 218.960 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 285.600 1099.000 286.160 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 1.000 995.120 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 796.000 706.160 799.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 20.160 1099.000 20.720 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 1.000 464.240 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 661.920 796.000 662.480 799.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 614.880 1099.000 615.440 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 221.760 1099.000 222.320 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 967.680 1.000 968.240 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1078.560 1.000 1079.120 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 154.560 4.000 155.120 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 920.640 1.000 921.200 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 141.120 1099.000 141.680 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 651.840 1099.000 652.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 1.000 54.320 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 1.000 393.680 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 796.000 296.240 799.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 796.000 286.160 799.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 675.360 4.000 675.920 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 1.000 218.960 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 1.000 857.360 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 688.800 796.000 689.360 799.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 796.000 477.680 799.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 796.000 114.800 799.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1014.720 1.000 1015.280 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 796.000 104.720 799.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 497.280 1099.000 497.840 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 796.000 507.920 799.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 77.280 1099.000 77.840 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 796.000 870.800 799.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 504.000 1099.000 504.560 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 362.880 4.000 363.440 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 413.280 1099.000 413.840 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 796.000 917.840 799.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 1.000 255.920 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 819.840 1.000 820.400 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1021.440 1.000 1022.000 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 120.960 1099.000 121.520 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1065.120 796.000 1065.680 799.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 53.760 4.000 54.320 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 305.760 1099.000 306.320 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 204.960 1099.000 205.520 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 524.160 1099.000 524.720 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 386.400 1099.000 386.960 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 796.000 158.480 799.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 756.000 4.000 756.560 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 1.000 702.800 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 1.000 840.560 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 1.000 134.960 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 117.600 4.000 118.160 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 796.000 215.600 799.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1031.520 1.000 1032.080 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 796.000 333.200 799.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 554.400 4.000 554.960 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 796.000 544.880 799.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 796.000 854.000 799.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 1.000 262.640 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 433.440 1099.000 434.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 1.000 850.640 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 796.000 343.280 799.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1.000 171.920 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 584.640 4.000 585.200 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 752.640 1099.000 753.200 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1092.000 796.000 1092.560 799.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 661.920 1099.000 662.480 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 796.000 561.680 799.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 624.960 1099.000 625.520 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 1.000 484.400 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 312.480 796.000 313.040 799.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1.000 27.440 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 1.000 7.280 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 796.000 279.440 799.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 1.000 491.120 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 409.920 4.000 410.480 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 520.800 4.000 521.360 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1068.480 1.000 1069.040 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 796.000 497.840 799.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 601.440 4.000 602.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 1.000 182.000 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.000 1.000 420.560 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 796.000 938.000 799.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 1.000 756.560 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.520 4.000 108.080 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 692.160 4.000 692.720 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 6.720 4.000 7.280 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 796.000 84.560 799.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 1.000 729.680 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 796.000 460.880 799.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 940.800 1.000 941.360 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 450.240 1099.000 450.800 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 510.720 4.000 511.280 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 339.360 1099.000 339.920 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 1.000 719.600 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 796.000 991.760 799.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1048.320 1.000 1048.880 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 796.000 716.240 799.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 1.000 877.520 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 463.680 4.000 464.240 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 1.000 118.160 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 322.560 1099.000 323.120 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.480 4.000 229.040 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 470.400 1099.000 470.960 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 1.000 235.760 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 1.000 904.400 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 796.000 423.920 799.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 964.320 796.000 964.880 799.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 577.920 1099.000 578.480 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 796.000 386.960 799.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 611.520 4.000 612.080 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 784.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 784.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 784.300 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 10.080 1099.000 10.640 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 796.000 323.120 799.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 174.720 1099.000 175.280 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 796.000 780.080 799.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 796.000 578.480 799.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 547.680 4.000 548.240 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 1.000 81.200 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 1.000 528.080 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 90.720 4.000 91.280 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 487.200 1099.000 487.760 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 1.000 602.000 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 527.520 4.000 528.080 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 147.840 1099.000 148.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 1.000 914.480 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 63.840 4.000 64.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1034.880 796.000 1035.440 799.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 1.000 538.160 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 766.080 1.000 766.640 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 67.200 1099.000 67.760 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 796.000 259.280 799.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 161.280 4.000 161.840 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 1.000 98.000 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 796.000 470.960 799.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 403.200 1099.000 403.760 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 762.720 1099.000 763.280 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 1.000 373.520 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 372.960 4.000 373.520 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 248.640 1099.000 249.200 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 1.000 739.760 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 796.000 880.880 799.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 1.000 712.880 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 235.200 4.000 235.760 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 1.000 44.240 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 1.000 951.440 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 104.160 1099.000 104.720 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 796.000 450.800 799.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 678.720 1099.000 679.280 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 729.120 4.000 729.680 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 796.000 3.920 799.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 766.080 4.000 766.640 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 1.000 34.160 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 198.240 4.000 198.800 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 349.440 1099.000 350.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 1.000 548.240 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 796.000 800.240 799.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 796.000 1028.720 799.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 796.000 205.520 799.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 1.000 145.040 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 446.880 4.000 447.440 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 796.000 1055.600 799.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 564.480 4.000 565.040 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 598.080 1099.000 598.640 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 157.920 1099.000 158.480 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 1.000 655.760 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 796.000 944.720 799.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 796.000 380.240 799.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 1.000 299.600 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 423.360 1099.000 423.920 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 1.000 776.720 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 131.040 1099.000 131.600 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 500.640 4.000 501.200 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 1.000 985.040 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 1.000 155.120 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 1.000 474.320 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 258.720 1099.000 259.280 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 900.480 796.000 901.040 799.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 698.880 1099.000 699.440 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 1.000 1005.200 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.520 4.000 192.080 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 396.480 1099.000 397.040 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1.000 17.360 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 725.760 1099.000 726.320 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 796.000 864.080 799.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1058.400 1.000 1058.960 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 796.000 837.200 799.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 262.080 4.000 262.640 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 299.040 4.000 299.600 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 1.000 638.960 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 1.000 749.840 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 456.960 4.000 457.520 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 796.000 20.720 799.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 796.000 413.840 799.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 309.120 4.000 309.680 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 1.000 198.800 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 1.000 71.120 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 796.000 642.320 799.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 796.000 434.000 799.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 1.000 521.360 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 806.400 796.000 806.960 799.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 110.880 1099.000 111.440 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 621.600 4.000 622.160 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 588.000 1099.000 588.560 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 1.000 208.880 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 1.000 363.440 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 80.640 4.000 81.200 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 551.040 1099.000 551.600 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 1.000 575.120 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 796.000 773.360 799.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 796.000 763.280 799.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 796.000 77.840 799.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 796.000 249.200 799.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 1.000 686.000 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 208.320 4.000 208.880 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 786.240 4.000 786.800 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1096.000 312.480 1099.000 313.040 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 1093.120 784.970 ;
      LAYER Metal2 ;
        RECT 0.140 795.700 3.060 796.000 ;
        RECT 4.220 795.700 13.140 796.000 ;
        RECT 14.300 795.700 19.860 796.000 ;
        RECT 21.020 795.700 29.940 796.000 ;
        RECT 31.100 795.700 40.020 796.000 ;
        RECT 41.180 795.700 50.100 796.000 ;
        RECT 51.260 795.700 56.820 796.000 ;
        RECT 57.980 795.700 66.900 796.000 ;
        RECT 68.060 795.700 76.980 796.000 ;
        RECT 78.140 795.700 83.700 796.000 ;
        RECT 84.860 795.700 93.780 796.000 ;
        RECT 94.940 795.700 103.860 796.000 ;
        RECT 105.020 795.700 113.940 796.000 ;
        RECT 115.100 795.700 120.660 796.000 ;
        RECT 121.820 795.700 130.740 796.000 ;
        RECT 131.900 795.700 140.820 796.000 ;
        RECT 141.980 795.700 147.540 796.000 ;
        RECT 148.700 795.700 157.620 796.000 ;
        RECT 158.780 795.700 167.700 796.000 ;
        RECT 168.860 795.700 177.780 796.000 ;
        RECT 178.940 795.700 184.500 796.000 ;
        RECT 185.660 795.700 194.580 796.000 ;
        RECT 195.740 795.700 204.660 796.000 ;
        RECT 205.820 795.700 214.740 796.000 ;
        RECT 215.900 795.700 221.460 796.000 ;
        RECT 222.620 795.700 231.540 796.000 ;
        RECT 232.700 795.700 241.620 796.000 ;
        RECT 242.780 795.700 248.340 796.000 ;
        RECT 249.500 795.700 258.420 796.000 ;
        RECT 259.580 795.700 268.500 796.000 ;
        RECT 269.660 795.700 278.580 796.000 ;
        RECT 279.740 795.700 285.300 796.000 ;
        RECT 286.460 795.700 295.380 796.000 ;
        RECT 296.540 795.700 305.460 796.000 ;
        RECT 306.620 795.700 312.180 796.000 ;
        RECT 313.340 795.700 322.260 796.000 ;
        RECT 323.420 795.700 332.340 796.000 ;
        RECT 333.500 795.700 342.420 796.000 ;
        RECT 343.580 795.700 349.140 796.000 ;
        RECT 350.300 795.700 359.220 796.000 ;
        RECT 360.380 795.700 369.300 796.000 ;
        RECT 370.460 795.700 379.380 796.000 ;
        RECT 380.540 795.700 386.100 796.000 ;
        RECT 387.260 795.700 396.180 796.000 ;
        RECT 397.340 795.700 406.260 796.000 ;
        RECT 407.420 795.700 412.980 796.000 ;
        RECT 414.140 795.700 423.060 796.000 ;
        RECT 424.220 795.700 433.140 796.000 ;
        RECT 434.300 795.700 443.220 796.000 ;
        RECT 444.380 795.700 449.940 796.000 ;
        RECT 451.100 795.700 460.020 796.000 ;
        RECT 461.180 795.700 470.100 796.000 ;
        RECT 471.260 795.700 476.820 796.000 ;
        RECT 477.980 795.700 486.900 796.000 ;
        RECT 488.060 795.700 496.980 796.000 ;
        RECT 498.140 795.700 507.060 796.000 ;
        RECT 508.220 795.700 513.780 796.000 ;
        RECT 514.940 795.700 523.860 796.000 ;
        RECT 525.020 795.700 533.940 796.000 ;
        RECT 535.100 795.700 544.020 796.000 ;
        RECT 545.180 795.700 550.740 796.000 ;
        RECT 551.900 795.700 560.820 796.000 ;
        RECT 561.980 795.700 570.900 796.000 ;
        RECT 572.060 795.700 577.620 796.000 ;
        RECT 578.780 795.700 587.700 796.000 ;
        RECT 588.860 795.700 597.780 796.000 ;
        RECT 598.940 795.700 607.860 796.000 ;
        RECT 609.020 795.700 614.580 796.000 ;
        RECT 615.740 795.700 624.660 796.000 ;
        RECT 625.820 795.700 634.740 796.000 ;
        RECT 635.900 795.700 641.460 796.000 ;
        RECT 642.620 795.700 651.540 796.000 ;
        RECT 652.700 795.700 661.620 796.000 ;
        RECT 662.780 795.700 671.700 796.000 ;
        RECT 672.860 795.700 678.420 796.000 ;
        RECT 679.580 795.700 688.500 796.000 ;
        RECT 689.660 795.700 698.580 796.000 ;
        RECT 699.740 795.700 705.300 796.000 ;
        RECT 706.460 795.700 715.380 796.000 ;
        RECT 716.540 795.700 725.460 796.000 ;
        RECT 726.620 795.700 735.540 796.000 ;
        RECT 736.700 795.700 742.260 796.000 ;
        RECT 743.420 795.700 752.340 796.000 ;
        RECT 753.500 795.700 762.420 796.000 ;
        RECT 763.580 795.700 772.500 796.000 ;
        RECT 773.660 795.700 779.220 796.000 ;
        RECT 780.380 795.700 789.300 796.000 ;
        RECT 790.460 795.700 799.380 796.000 ;
        RECT 800.540 795.700 806.100 796.000 ;
        RECT 807.260 795.700 816.180 796.000 ;
        RECT 817.340 795.700 826.260 796.000 ;
        RECT 827.420 795.700 836.340 796.000 ;
        RECT 837.500 795.700 843.060 796.000 ;
        RECT 844.220 795.700 853.140 796.000 ;
        RECT 854.300 795.700 863.220 796.000 ;
        RECT 864.380 795.700 869.940 796.000 ;
        RECT 871.100 795.700 880.020 796.000 ;
        RECT 881.180 795.700 890.100 796.000 ;
        RECT 891.260 795.700 900.180 796.000 ;
        RECT 901.340 795.700 906.900 796.000 ;
        RECT 908.060 795.700 916.980 796.000 ;
        RECT 918.140 795.700 927.060 796.000 ;
        RECT 928.220 795.700 937.140 796.000 ;
        RECT 938.300 795.700 943.860 796.000 ;
        RECT 945.020 795.700 953.940 796.000 ;
        RECT 955.100 795.700 964.020 796.000 ;
        RECT 965.180 795.700 970.740 796.000 ;
        RECT 971.900 795.700 980.820 796.000 ;
        RECT 981.980 795.700 990.900 796.000 ;
        RECT 992.060 795.700 1000.980 796.000 ;
        RECT 1002.140 795.700 1007.700 796.000 ;
        RECT 1008.860 795.700 1017.780 796.000 ;
        RECT 1018.940 795.700 1027.860 796.000 ;
        RECT 1029.020 795.700 1034.580 796.000 ;
        RECT 1035.740 795.700 1044.660 796.000 ;
        RECT 1045.820 795.700 1054.740 796.000 ;
        RECT 1055.900 795.700 1064.820 796.000 ;
        RECT 1065.980 795.700 1071.540 796.000 ;
        RECT 1072.700 795.700 1081.620 796.000 ;
        RECT 1082.780 795.700 1090.740 796.000 ;
        RECT 0.140 4.300 1090.740 795.700 ;
        RECT 0.860 4.000 6.420 4.300 ;
        RECT 7.580 4.000 16.500 4.300 ;
        RECT 17.660 4.000 26.580 4.300 ;
        RECT 27.740 4.000 33.300 4.300 ;
        RECT 34.460 4.000 43.380 4.300 ;
        RECT 44.540 4.000 53.460 4.300 ;
        RECT 54.620 4.000 63.540 4.300 ;
        RECT 64.700 4.000 70.260 4.300 ;
        RECT 71.420 4.000 80.340 4.300 ;
        RECT 81.500 4.000 90.420 4.300 ;
        RECT 91.580 4.000 97.140 4.300 ;
        RECT 98.300 4.000 107.220 4.300 ;
        RECT 108.380 4.000 117.300 4.300 ;
        RECT 118.460 4.000 127.380 4.300 ;
        RECT 128.540 4.000 134.100 4.300 ;
        RECT 135.260 4.000 144.180 4.300 ;
        RECT 145.340 4.000 154.260 4.300 ;
        RECT 155.420 4.000 160.980 4.300 ;
        RECT 162.140 4.000 171.060 4.300 ;
        RECT 172.220 4.000 181.140 4.300 ;
        RECT 182.300 4.000 191.220 4.300 ;
        RECT 192.380 4.000 197.940 4.300 ;
        RECT 199.100 4.000 208.020 4.300 ;
        RECT 209.180 4.000 218.100 4.300 ;
        RECT 219.260 4.000 228.180 4.300 ;
        RECT 229.340 4.000 234.900 4.300 ;
        RECT 236.060 4.000 244.980 4.300 ;
        RECT 246.140 4.000 255.060 4.300 ;
        RECT 256.220 4.000 261.780 4.300 ;
        RECT 262.940 4.000 271.860 4.300 ;
        RECT 273.020 4.000 281.940 4.300 ;
        RECT 283.100 4.000 292.020 4.300 ;
        RECT 293.180 4.000 298.740 4.300 ;
        RECT 299.900 4.000 308.820 4.300 ;
        RECT 309.980 4.000 318.900 4.300 ;
        RECT 320.060 4.000 325.620 4.300 ;
        RECT 326.780 4.000 335.700 4.300 ;
        RECT 336.860 4.000 345.780 4.300 ;
        RECT 346.940 4.000 355.860 4.300 ;
        RECT 357.020 4.000 362.580 4.300 ;
        RECT 363.740 4.000 372.660 4.300 ;
        RECT 373.820 4.000 382.740 4.300 ;
        RECT 383.900 4.000 392.820 4.300 ;
        RECT 393.980 4.000 399.540 4.300 ;
        RECT 400.700 4.000 409.620 4.300 ;
        RECT 410.780 4.000 419.700 4.300 ;
        RECT 420.860 4.000 426.420 4.300 ;
        RECT 427.580 4.000 436.500 4.300 ;
        RECT 437.660 4.000 446.580 4.300 ;
        RECT 447.740 4.000 456.660 4.300 ;
        RECT 457.820 4.000 463.380 4.300 ;
        RECT 464.540 4.000 473.460 4.300 ;
        RECT 474.620 4.000 483.540 4.300 ;
        RECT 484.700 4.000 490.260 4.300 ;
        RECT 491.420 4.000 500.340 4.300 ;
        RECT 501.500 4.000 510.420 4.300 ;
        RECT 511.580 4.000 520.500 4.300 ;
        RECT 521.660 4.000 527.220 4.300 ;
        RECT 528.380 4.000 537.300 4.300 ;
        RECT 538.460 4.000 547.380 4.300 ;
        RECT 548.540 4.000 554.100 4.300 ;
        RECT 555.260 4.000 564.180 4.300 ;
        RECT 565.340 4.000 574.260 4.300 ;
        RECT 575.420 4.000 584.340 4.300 ;
        RECT 585.500 4.000 591.060 4.300 ;
        RECT 592.220 4.000 601.140 4.300 ;
        RECT 602.300 4.000 611.220 4.300 ;
        RECT 612.380 4.000 621.300 4.300 ;
        RECT 622.460 4.000 628.020 4.300 ;
        RECT 629.180 4.000 638.100 4.300 ;
        RECT 639.260 4.000 648.180 4.300 ;
        RECT 649.340 4.000 654.900 4.300 ;
        RECT 656.060 4.000 664.980 4.300 ;
        RECT 666.140 4.000 675.060 4.300 ;
        RECT 676.220 4.000 685.140 4.300 ;
        RECT 686.300 4.000 691.860 4.300 ;
        RECT 693.020 4.000 701.940 4.300 ;
        RECT 703.100 4.000 712.020 4.300 ;
        RECT 713.180 4.000 718.740 4.300 ;
        RECT 719.900 4.000 728.820 4.300 ;
        RECT 729.980 4.000 738.900 4.300 ;
        RECT 740.060 4.000 748.980 4.300 ;
        RECT 750.140 4.000 755.700 4.300 ;
        RECT 756.860 4.000 765.780 4.300 ;
        RECT 766.940 4.000 775.860 4.300 ;
        RECT 777.020 4.000 785.940 4.300 ;
        RECT 787.100 4.000 792.660 4.300 ;
        RECT 793.820 4.000 802.740 4.300 ;
        RECT 803.900 4.000 812.820 4.300 ;
        RECT 813.980 4.000 819.540 4.300 ;
        RECT 820.700 4.000 829.620 4.300 ;
        RECT 830.780 4.000 839.700 4.300 ;
        RECT 840.860 4.000 849.780 4.300 ;
        RECT 850.940 4.000 856.500 4.300 ;
        RECT 857.660 4.000 866.580 4.300 ;
        RECT 867.740 4.000 876.660 4.300 ;
        RECT 877.820 4.000 883.380 4.300 ;
        RECT 884.540 4.000 893.460 4.300 ;
        RECT 894.620 4.000 903.540 4.300 ;
        RECT 904.700 4.000 913.620 4.300 ;
        RECT 914.780 4.000 920.340 4.300 ;
        RECT 921.500 4.000 930.420 4.300 ;
        RECT 931.580 4.000 940.500 4.300 ;
        RECT 941.660 4.000 950.580 4.300 ;
        RECT 951.740 4.000 957.300 4.300 ;
        RECT 958.460 4.000 967.380 4.300 ;
        RECT 968.540 4.000 977.460 4.300 ;
        RECT 978.620 4.000 984.180 4.300 ;
        RECT 985.340 4.000 994.260 4.300 ;
        RECT 995.420 4.000 1004.340 4.300 ;
        RECT 1005.500 4.000 1014.420 4.300 ;
        RECT 1015.580 4.000 1021.140 4.300 ;
        RECT 1022.300 4.000 1031.220 4.300 ;
        RECT 1032.380 4.000 1041.300 4.300 ;
        RECT 1042.460 4.000 1048.020 4.300 ;
        RECT 1049.180 4.000 1058.100 4.300 ;
        RECT 1059.260 4.000 1068.180 4.300 ;
        RECT 1069.340 4.000 1078.260 4.300 ;
        RECT 1079.420 4.000 1084.980 4.300 ;
        RECT 1086.140 4.000 1090.740 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 780.380 1099.700 784.140 ;
        RECT 0.090 779.220 1095.700 780.380 ;
        RECT 1099.300 779.220 1099.700 780.380 ;
        RECT 0.090 777.020 1099.700 779.220 ;
        RECT 0.090 775.860 0.700 777.020 ;
        RECT 4.300 775.860 1099.700 777.020 ;
        RECT 0.090 770.300 1099.700 775.860 ;
        RECT 0.090 769.140 1095.700 770.300 ;
        RECT 1099.300 769.140 1099.700 770.300 ;
        RECT 0.090 766.940 1099.700 769.140 ;
        RECT 0.090 765.780 0.700 766.940 ;
        RECT 4.300 765.780 1099.700 766.940 ;
        RECT 0.090 763.580 1099.700 765.780 ;
        RECT 0.090 762.420 1095.700 763.580 ;
        RECT 1099.300 762.420 1099.700 763.580 ;
        RECT 0.090 756.860 1099.700 762.420 ;
        RECT 0.090 755.700 0.700 756.860 ;
        RECT 4.300 755.700 1099.700 756.860 ;
        RECT 0.090 753.500 1099.700 755.700 ;
        RECT 0.090 752.340 1095.700 753.500 ;
        RECT 1099.300 752.340 1099.700 753.500 ;
        RECT 0.090 750.140 1099.700 752.340 ;
        RECT 0.090 748.980 0.700 750.140 ;
        RECT 4.300 748.980 1099.700 750.140 ;
        RECT 0.090 743.420 1099.700 748.980 ;
        RECT 0.090 742.260 1095.700 743.420 ;
        RECT 1099.300 742.260 1099.700 743.420 ;
        RECT 0.090 740.060 1099.700 742.260 ;
        RECT 0.090 738.900 0.700 740.060 ;
        RECT 4.300 738.900 1099.700 740.060 ;
        RECT 0.090 733.340 1099.700 738.900 ;
        RECT 0.090 732.180 1095.700 733.340 ;
        RECT 1099.300 732.180 1099.700 733.340 ;
        RECT 0.090 729.980 1099.700 732.180 ;
        RECT 0.090 728.820 0.700 729.980 ;
        RECT 4.300 728.820 1099.700 729.980 ;
        RECT 0.090 726.620 1099.700 728.820 ;
        RECT 0.090 725.460 1095.700 726.620 ;
        RECT 1099.300 725.460 1099.700 726.620 ;
        RECT 0.090 719.900 1099.700 725.460 ;
        RECT 0.090 718.740 0.700 719.900 ;
        RECT 4.300 718.740 1099.700 719.900 ;
        RECT 0.090 716.540 1099.700 718.740 ;
        RECT 0.090 715.380 1095.700 716.540 ;
        RECT 1099.300 715.380 1099.700 716.540 ;
        RECT 0.090 713.180 1099.700 715.380 ;
        RECT 0.090 712.020 0.700 713.180 ;
        RECT 4.300 712.020 1099.700 713.180 ;
        RECT 0.090 706.460 1099.700 712.020 ;
        RECT 0.090 705.300 1095.700 706.460 ;
        RECT 1099.300 705.300 1099.700 706.460 ;
        RECT 0.090 703.100 1099.700 705.300 ;
        RECT 0.090 701.940 0.700 703.100 ;
        RECT 4.300 701.940 1099.700 703.100 ;
        RECT 0.090 699.740 1099.700 701.940 ;
        RECT 0.090 698.580 1095.700 699.740 ;
        RECT 1099.300 698.580 1099.700 699.740 ;
        RECT 0.090 693.020 1099.700 698.580 ;
        RECT 0.090 691.860 0.700 693.020 ;
        RECT 4.300 691.860 1099.700 693.020 ;
        RECT 0.090 689.660 1099.700 691.860 ;
        RECT 0.090 688.500 1095.700 689.660 ;
        RECT 1099.300 688.500 1099.700 689.660 ;
        RECT 0.090 686.300 1099.700 688.500 ;
        RECT 0.090 685.140 0.700 686.300 ;
        RECT 4.300 685.140 1099.700 686.300 ;
        RECT 0.090 679.580 1099.700 685.140 ;
        RECT 0.090 678.420 1095.700 679.580 ;
        RECT 1099.300 678.420 1099.700 679.580 ;
        RECT 0.090 676.220 1099.700 678.420 ;
        RECT 0.090 675.060 0.700 676.220 ;
        RECT 4.300 675.060 1099.700 676.220 ;
        RECT 0.090 669.500 1099.700 675.060 ;
        RECT 0.090 668.340 1095.700 669.500 ;
        RECT 1099.300 668.340 1099.700 669.500 ;
        RECT 0.090 666.140 1099.700 668.340 ;
        RECT 0.090 664.980 0.700 666.140 ;
        RECT 4.300 664.980 1099.700 666.140 ;
        RECT 0.090 662.780 1099.700 664.980 ;
        RECT 0.090 661.620 1095.700 662.780 ;
        RECT 1099.300 661.620 1099.700 662.780 ;
        RECT 0.090 656.060 1099.700 661.620 ;
        RECT 0.090 654.900 0.700 656.060 ;
        RECT 4.300 654.900 1099.700 656.060 ;
        RECT 0.090 652.700 1099.700 654.900 ;
        RECT 0.090 651.540 1095.700 652.700 ;
        RECT 1099.300 651.540 1099.700 652.700 ;
        RECT 0.090 649.340 1099.700 651.540 ;
        RECT 0.090 648.180 0.700 649.340 ;
        RECT 4.300 648.180 1099.700 649.340 ;
        RECT 0.090 642.620 1099.700 648.180 ;
        RECT 0.090 641.460 1095.700 642.620 ;
        RECT 1099.300 641.460 1099.700 642.620 ;
        RECT 0.090 639.260 1099.700 641.460 ;
        RECT 0.090 638.100 0.700 639.260 ;
        RECT 4.300 638.100 1099.700 639.260 ;
        RECT 0.090 635.900 1099.700 638.100 ;
        RECT 0.090 634.740 1095.700 635.900 ;
        RECT 1099.300 634.740 1099.700 635.900 ;
        RECT 0.090 629.180 1099.700 634.740 ;
        RECT 0.090 628.020 0.700 629.180 ;
        RECT 4.300 628.020 1099.700 629.180 ;
        RECT 0.090 625.820 1099.700 628.020 ;
        RECT 0.090 624.660 1095.700 625.820 ;
        RECT 1099.300 624.660 1099.700 625.820 ;
        RECT 0.090 622.460 1099.700 624.660 ;
        RECT 0.090 621.300 0.700 622.460 ;
        RECT 4.300 621.300 1099.700 622.460 ;
        RECT 0.090 615.740 1099.700 621.300 ;
        RECT 0.090 614.580 1095.700 615.740 ;
        RECT 1099.300 614.580 1099.700 615.740 ;
        RECT 0.090 612.380 1099.700 614.580 ;
        RECT 0.090 611.220 0.700 612.380 ;
        RECT 4.300 611.220 1099.700 612.380 ;
        RECT 0.090 605.660 1099.700 611.220 ;
        RECT 0.090 604.500 1095.700 605.660 ;
        RECT 1099.300 604.500 1099.700 605.660 ;
        RECT 0.090 602.300 1099.700 604.500 ;
        RECT 0.090 601.140 0.700 602.300 ;
        RECT 4.300 601.140 1099.700 602.300 ;
        RECT 0.090 598.940 1099.700 601.140 ;
        RECT 0.090 597.780 1095.700 598.940 ;
        RECT 1099.300 597.780 1099.700 598.940 ;
        RECT 0.090 592.220 1099.700 597.780 ;
        RECT 0.090 591.060 0.700 592.220 ;
        RECT 4.300 591.060 1099.700 592.220 ;
        RECT 0.090 588.860 1099.700 591.060 ;
        RECT 0.090 587.700 1095.700 588.860 ;
        RECT 1099.300 587.700 1099.700 588.860 ;
        RECT 0.090 585.500 1099.700 587.700 ;
        RECT 0.090 584.340 0.700 585.500 ;
        RECT 4.300 584.340 1099.700 585.500 ;
        RECT 0.090 578.780 1099.700 584.340 ;
        RECT 0.090 577.620 1095.700 578.780 ;
        RECT 1099.300 577.620 1099.700 578.780 ;
        RECT 0.090 575.420 1099.700 577.620 ;
        RECT 0.090 574.260 0.700 575.420 ;
        RECT 4.300 574.260 1099.700 575.420 ;
        RECT 0.090 568.700 1099.700 574.260 ;
        RECT 0.090 567.540 1095.700 568.700 ;
        RECT 1099.300 567.540 1099.700 568.700 ;
        RECT 0.090 565.340 1099.700 567.540 ;
        RECT 0.090 564.180 0.700 565.340 ;
        RECT 4.300 564.180 1099.700 565.340 ;
        RECT 0.090 561.980 1099.700 564.180 ;
        RECT 0.090 560.820 1095.700 561.980 ;
        RECT 1099.300 560.820 1099.700 561.980 ;
        RECT 0.090 555.260 1099.700 560.820 ;
        RECT 0.090 554.100 0.700 555.260 ;
        RECT 4.300 554.100 1099.700 555.260 ;
        RECT 0.090 551.900 1099.700 554.100 ;
        RECT 0.090 550.740 1095.700 551.900 ;
        RECT 1099.300 550.740 1099.700 551.900 ;
        RECT 0.090 548.540 1099.700 550.740 ;
        RECT 0.090 547.380 0.700 548.540 ;
        RECT 4.300 547.380 1099.700 548.540 ;
        RECT 0.090 541.820 1099.700 547.380 ;
        RECT 0.090 540.660 1095.700 541.820 ;
        RECT 1099.300 540.660 1099.700 541.820 ;
        RECT 0.090 538.460 1099.700 540.660 ;
        RECT 0.090 537.300 0.700 538.460 ;
        RECT 4.300 537.300 1099.700 538.460 ;
        RECT 0.090 535.100 1099.700 537.300 ;
        RECT 0.090 533.940 1095.700 535.100 ;
        RECT 1099.300 533.940 1099.700 535.100 ;
        RECT 0.090 528.380 1099.700 533.940 ;
        RECT 0.090 527.220 0.700 528.380 ;
        RECT 4.300 527.220 1099.700 528.380 ;
        RECT 0.090 525.020 1099.700 527.220 ;
        RECT 0.090 523.860 1095.700 525.020 ;
        RECT 1099.300 523.860 1099.700 525.020 ;
        RECT 0.090 521.660 1099.700 523.860 ;
        RECT 0.090 520.500 0.700 521.660 ;
        RECT 4.300 520.500 1099.700 521.660 ;
        RECT 0.090 514.940 1099.700 520.500 ;
        RECT 0.090 513.780 1095.700 514.940 ;
        RECT 1099.300 513.780 1099.700 514.940 ;
        RECT 0.090 511.580 1099.700 513.780 ;
        RECT 0.090 510.420 0.700 511.580 ;
        RECT 4.300 510.420 1099.700 511.580 ;
        RECT 0.090 504.860 1099.700 510.420 ;
        RECT 0.090 503.700 1095.700 504.860 ;
        RECT 1099.300 503.700 1099.700 504.860 ;
        RECT 0.090 501.500 1099.700 503.700 ;
        RECT 0.090 500.340 0.700 501.500 ;
        RECT 4.300 500.340 1099.700 501.500 ;
        RECT 0.090 498.140 1099.700 500.340 ;
        RECT 0.090 496.980 1095.700 498.140 ;
        RECT 1099.300 496.980 1099.700 498.140 ;
        RECT 0.090 491.420 1099.700 496.980 ;
        RECT 0.090 490.260 0.700 491.420 ;
        RECT 4.300 490.260 1099.700 491.420 ;
        RECT 0.090 488.060 1099.700 490.260 ;
        RECT 0.090 486.900 1095.700 488.060 ;
        RECT 1099.300 486.900 1099.700 488.060 ;
        RECT 0.090 484.700 1099.700 486.900 ;
        RECT 0.090 483.540 0.700 484.700 ;
        RECT 4.300 483.540 1099.700 484.700 ;
        RECT 0.090 477.980 1099.700 483.540 ;
        RECT 0.090 476.820 1095.700 477.980 ;
        RECT 1099.300 476.820 1099.700 477.980 ;
        RECT 0.090 474.620 1099.700 476.820 ;
        RECT 0.090 473.460 0.700 474.620 ;
        RECT 4.300 473.460 1099.700 474.620 ;
        RECT 0.090 471.260 1099.700 473.460 ;
        RECT 0.090 470.100 1095.700 471.260 ;
        RECT 1099.300 470.100 1099.700 471.260 ;
        RECT 0.090 464.540 1099.700 470.100 ;
        RECT 0.090 463.380 0.700 464.540 ;
        RECT 4.300 463.380 1099.700 464.540 ;
        RECT 0.090 461.180 1099.700 463.380 ;
        RECT 0.090 460.020 1095.700 461.180 ;
        RECT 1099.300 460.020 1099.700 461.180 ;
        RECT 0.090 457.820 1099.700 460.020 ;
        RECT 0.090 456.660 0.700 457.820 ;
        RECT 4.300 456.660 1099.700 457.820 ;
        RECT 0.090 451.100 1099.700 456.660 ;
        RECT 0.090 449.940 1095.700 451.100 ;
        RECT 1099.300 449.940 1099.700 451.100 ;
        RECT 0.090 447.740 1099.700 449.940 ;
        RECT 0.090 446.580 0.700 447.740 ;
        RECT 4.300 446.580 1099.700 447.740 ;
        RECT 0.090 441.020 1099.700 446.580 ;
        RECT 0.090 439.860 1095.700 441.020 ;
        RECT 1099.300 439.860 1099.700 441.020 ;
        RECT 0.090 437.660 1099.700 439.860 ;
        RECT 0.090 436.500 0.700 437.660 ;
        RECT 4.300 436.500 1099.700 437.660 ;
        RECT 0.090 434.300 1099.700 436.500 ;
        RECT 0.090 433.140 1095.700 434.300 ;
        RECT 1099.300 433.140 1099.700 434.300 ;
        RECT 0.090 427.580 1099.700 433.140 ;
        RECT 0.090 426.420 0.700 427.580 ;
        RECT 4.300 426.420 1099.700 427.580 ;
        RECT 0.090 424.220 1099.700 426.420 ;
        RECT 0.090 423.060 1095.700 424.220 ;
        RECT 1099.300 423.060 1099.700 424.220 ;
        RECT 0.090 420.860 1099.700 423.060 ;
        RECT 0.090 419.700 0.700 420.860 ;
        RECT 4.300 419.700 1099.700 420.860 ;
        RECT 0.090 414.140 1099.700 419.700 ;
        RECT 0.090 412.980 1095.700 414.140 ;
        RECT 1099.300 412.980 1099.700 414.140 ;
        RECT 0.090 410.780 1099.700 412.980 ;
        RECT 0.090 409.620 0.700 410.780 ;
        RECT 4.300 409.620 1099.700 410.780 ;
        RECT 0.090 404.060 1099.700 409.620 ;
        RECT 0.090 402.900 1095.700 404.060 ;
        RECT 1099.300 402.900 1099.700 404.060 ;
        RECT 0.090 400.700 1099.700 402.900 ;
        RECT 0.090 399.540 0.700 400.700 ;
        RECT 4.300 399.540 1099.700 400.700 ;
        RECT 0.090 397.340 1099.700 399.540 ;
        RECT 0.090 396.180 1095.700 397.340 ;
        RECT 1099.300 396.180 1099.700 397.340 ;
        RECT 0.090 393.980 1099.700 396.180 ;
        RECT 0.090 392.820 0.700 393.980 ;
        RECT 4.300 392.820 1099.700 393.980 ;
        RECT 0.090 387.260 1099.700 392.820 ;
        RECT 0.090 386.100 1095.700 387.260 ;
        RECT 1099.300 386.100 1099.700 387.260 ;
        RECT 0.090 383.900 1099.700 386.100 ;
        RECT 0.090 382.740 0.700 383.900 ;
        RECT 4.300 382.740 1099.700 383.900 ;
        RECT 0.090 377.180 1099.700 382.740 ;
        RECT 0.090 376.020 1095.700 377.180 ;
        RECT 1099.300 376.020 1099.700 377.180 ;
        RECT 0.090 373.820 1099.700 376.020 ;
        RECT 0.090 372.660 0.700 373.820 ;
        RECT 4.300 372.660 1099.700 373.820 ;
        RECT 0.090 370.460 1099.700 372.660 ;
        RECT 0.090 369.300 1095.700 370.460 ;
        RECT 1099.300 369.300 1099.700 370.460 ;
        RECT 0.090 363.740 1099.700 369.300 ;
        RECT 0.090 362.580 0.700 363.740 ;
        RECT 4.300 362.580 1099.700 363.740 ;
        RECT 0.090 360.380 1099.700 362.580 ;
        RECT 0.090 359.220 1095.700 360.380 ;
        RECT 1099.300 359.220 1099.700 360.380 ;
        RECT 0.090 357.020 1099.700 359.220 ;
        RECT 0.090 355.860 0.700 357.020 ;
        RECT 4.300 355.860 1099.700 357.020 ;
        RECT 0.090 350.300 1099.700 355.860 ;
        RECT 0.090 349.140 1095.700 350.300 ;
        RECT 1099.300 349.140 1099.700 350.300 ;
        RECT 0.090 346.940 1099.700 349.140 ;
        RECT 0.090 345.780 0.700 346.940 ;
        RECT 4.300 345.780 1099.700 346.940 ;
        RECT 0.090 340.220 1099.700 345.780 ;
        RECT 0.090 339.060 1095.700 340.220 ;
        RECT 1099.300 339.060 1099.700 340.220 ;
        RECT 0.090 336.860 1099.700 339.060 ;
        RECT 0.090 335.700 0.700 336.860 ;
        RECT 4.300 335.700 1099.700 336.860 ;
        RECT 0.090 333.500 1099.700 335.700 ;
        RECT 0.090 332.340 1095.700 333.500 ;
        RECT 1099.300 332.340 1099.700 333.500 ;
        RECT 0.090 326.780 1099.700 332.340 ;
        RECT 0.090 325.620 0.700 326.780 ;
        RECT 4.300 325.620 1099.700 326.780 ;
        RECT 0.090 323.420 1099.700 325.620 ;
        RECT 0.090 322.260 1095.700 323.420 ;
        RECT 1099.300 322.260 1099.700 323.420 ;
        RECT 0.090 320.060 1099.700 322.260 ;
        RECT 0.090 318.900 0.700 320.060 ;
        RECT 4.300 318.900 1099.700 320.060 ;
        RECT 0.090 313.340 1099.700 318.900 ;
        RECT 0.090 312.180 1095.700 313.340 ;
        RECT 1099.300 312.180 1099.700 313.340 ;
        RECT 0.090 309.980 1099.700 312.180 ;
        RECT 0.090 308.820 0.700 309.980 ;
        RECT 4.300 308.820 1099.700 309.980 ;
        RECT 0.090 306.620 1099.700 308.820 ;
        RECT 0.090 305.460 1095.700 306.620 ;
        RECT 1099.300 305.460 1099.700 306.620 ;
        RECT 0.090 299.900 1099.700 305.460 ;
        RECT 0.090 298.740 0.700 299.900 ;
        RECT 4.300 298.740 1099.700 299.900 ;
        RECT 0.090 296.540 1099.700 298.740 ;
        RECT 0.090 295.380 1095.700 296.540 ;
        RECT 1099.300 295.380 1099.700 296.540 ;
        RECT 0.090 293.180 1099.700 295.380 ;
        RECT 0.090 292.020 0.700 293.180 ;
        RECT 4.300 292.020 1099.700 293.180 ;
        RECT 0.090 286.460 1099.700 292.020 ;
        RECT 0.090 285.300 1095.700 286.460 ;
        RECT 1099.300 285.300 1099.700 286.460 ;
        RECT 0.090 283.100 1099.700 285.300 ;
        RECT 0.090 281.940 0.700 283.100 ;
        RECT 4.300 281.940 1099.700 283.100 ;
        RECT 0.090 276.380 1099.700 281.940 ;
        RECT 0.090 275.220 1095.700 276.380 ;
        RECT 1099.300 275.220 1099.700 276.380 ;
        RECT 0.090 273.020 1099.700 275.220 ;
        RECT 0.090 271.860 0.700 273.020 ;
        RECT 4.300 271.860 1099.700 273.020 ;
        RECT 0.090 269.660 1099.700 271.860 ;
        RECT 0.090 268.500 1095.700 269.660 ;
        RECT 1099.300 268.500 1099.700 269.660 ;
        RECT 0.090 262.940 1099.700 268.500 ;
        RECT 0.090 261.780 0.700 262.940 ;
        RECT 4.300 261.780 1099.700 262.940 ;
        RECT 0.090 259.580 1099.700 261.780 ;
        RECT 0.090 258.420 1095.700 259.580 ;
        RECT 1099.300 258.420 1099.700 259.580 ;
        RECT 0.090 256.220 1099.700 258.420 ;
        RECT 0.090 255.060 0.700 256.220 ;
        RECT 4.300 255.060 1099.700 256.220 ;
        RECT 0.090 249.500 1099.700 255.060 ;
        RECT 0.090 248.340 1095.700 249.500 ;
        RECT 1099.300 248.340 1099.700 249.500 ;
        RECT 0.090 246.140 1099.700 248.340 ;
        RECT 0.090 244.980 0.700 246.140 ;
        RECT 4.300 244.980 1099.700 246.140 ;
        RECT 0.090 242.780 1099.700 244.980 ;
        RECT 0.090 241.620 1095.700 242.780 ;
        RECT 1099.300 241.620 1099.700 242.780 ;
        RECT 0.090 236.060 1099.700 241.620 ;
        RECT 0.090 234.900 0.700 236.060 ;
        RECT 4.300 234.900 1099.700 236.060 ;
        RECT 0.090 232.700 1099.700 234.900 ;
        RECT 0.090 231.540 1095.700 232.700 ;
        RECT 1099.300 231.540 1099.700 232.700 ;
        RECT 0.090 229.340 1099.700 231.540 ;
        RECT 0.090 228.180 0.700 229.340 ;
        RECT 4.300 228.180 1099.700 229.340 ;
        RECT 0.090 222.620 1099.700 228.180 ;
        RECT 0.090 221.460 1095.700 222.620 ;
        RECT 1099.300 221.460 1099.700 222.620 ;
        RECT 0.090 219.260 1099.700 221.460 ;
        RECT 0.090 218.100 0.700 219.260 ;
        RECT 4.300 218.100 1099.700 219.260 ;
        RECT 0.090 212.540 1099.700 218.100 ;
        RECT 0.090 211.380 1095.700 212.540 ;
        RECT 1099.300 211.380 1099.700 212.540 ;
        RECT 0.090 209.180 1099.700 211.380 ;
        RECT 0.090 208.020 0.700 209.180 ;
        RECT 4.300 208.020 1099.700 209.180 ;
        RECT 0.090 205.820 1099.700 208.020 ;
        RECT 0.090 204.660 1095.700 205.820 ;
        RECT 1099.300 204.660 1099.700 205.820 ;
        RECT 0.090 199.100 1099.700 204.660 ;
        RECT 0.090 197.940 0.700 199.100 ;
        RECT 4.300 197.940 1099.700 199.100 ;
        RECT 0.090 195.740 1099.700 197.940 ;
        RECT 0.090 194.580 1095.700 195.740 ;
        RECT 1099.300 194.580 1099.700 195.740 ;
        RECT 0.090 192.380 1099.700 194.580 ;
        RECT 0.090 191.220 0.700 192.380 ;
        RECT 4.300 191.220 1099.700 192.380 ;
        RECT 0.090 185.660 1099.700 191.220 ;
        RECT 0.090 184.500 1095.700 185.660 ;
        RECT 1099.300 184.500 1099.700 185.660 ;
        RECT 0.090 182.300 1099.700 184.500 ;
        RECT 0.090 181.140 0.700 182.300 ;
        RECT 4.300 181.140 1099.700 182.300 ;
        RECT 0.090 175.580 1099.700 181.140 ;
        RECT 0.090 174.420 1095.700 175.580 ;
        RECT 1099.300 174.420 1099.700 175.580 ;
        RECT 0.090 172.220 1099.700 174.420 ;
        RECT 0.090 171.060 0.700 172.220 ;
        RECT 4.300 171.060 1099.700 172.220 ;
        RECT 0.090 168.860 1099.700 171.060 ;
        RECT 0.090 167.700 1095.700 168.860 ;
        RECT 1099.300 167.700 1099.700 168.860 ;
        RECT 0.090 162.140 1099.700 167.700 ;
        RECT 0.090 160.980 0.700 162.140 ;
        RECT 4.300 160.980 1099.700 162.140 ;
        RECT 0.090 158.780 1099.700 160.980 ;
        RECT 0.090 157.620 1095.700 158.780 ;
        RECT 1099.300 157.620 1099.700 158.780 ;
        RECT 0.090 155.420 1099.700 157.620 ;
        RECT 0.090 154.260 0.700 155.420 ;
        RECT 4.300 154.260 1099.700 155.420 ;
        RECT 0.090 148.700 1099.700 154.260 ;
        RECT 0.090 147.540 1095.700 148.700 ;
        RECT 1099.300 147.540 1099.700 148.700 ;
        RECT 0.090 145.340 1099.700 147.540 ;
        RECT 0.090 144.180 0.700 145.340 ;
        RECT 4.300 144.180 1099.700 145.340 ;
        RECT 0.090 141.980 1099.700 144.180 ;
        RECT 0.090 140.820 1095.700 141.980 ;
        RECT 1099.300 140.820 1099.700 141.980 ;
        RECT 0.090 135.260 1099.700 140.820 ;
        RECT 0.090 134.100 0.700 135.260 ;
        RECT 4.300 134.100 1099.700 135.260 ;
        RECT 0.090 131.900 1099.700 134.100 ;
        RECT 0.090 130.740 1095.700 131.900 ;
        RECT 1099.300 130.740 1099.700 131.900 ;
        RECT 0.090 128.540 1099.700 130.740 ;
        RECT 0.090 127.380 0.700 128.540 ;
        RECT 4.300 127.380 1099.700 128.540 ;
        RECT 0.090 121.820 1099.700 127.380 ;
        RECT 0.090 120.660 1095.700 121.820 ;
        RECT 1099.300 120.660 1099.700 121.820 ;
        RECT 0.090 118.460 1099.700 120.660 ;
        RECT 0.090 117.300 0.700 118.460 ;
        RECT 4.300 117.300 1099.700 118.460 ;
        RECT 0.090 111.740 1099.700 117.300 ;
        RECT 0.090 110.580 1095.700 111.740 ;
        RECT 1099.300 110.580 1099.700 111.740 ;
        RECT 0.090 108.380 1099.700 110.580 ;
        RECT 0.090 107.220 0.700 108.380 ;
        RECT 4.300 107.220 1099.700 108.380 ;
        RECT 0.090 105.020 1099.700 107.220 ;
        RECT 0.090 103.860 1095.700 105.020 ;
        RECT 1099.300 103.860 1099.700 105.020 ;
        RECT 0.090 98.300 1099.700 103.860 ;
        RECT 0.090 97.140 0.700 98.300 ;
        RECT 4.300 97.140 1099.700 98.300 ;
        RECT 0.090 94.940 1099.700 97.140 ;
        RECT 0.090 93.780 1095.700 94.940 ;
        RECT 1099.300 93.780 1099.700 94.940 ;
        RECT 0.090 91.580 1099.700 93.780 ;
        RECT 0.090 90.420 0.700 91.580 ;
        RECT 4.300 90.420 1099.700 91.580 ;
        RECT 0.090 84.860 1099.700 90.420 ;
        RECT 0.090 83.700 1095.700 84.860 ;
        RECT 1099.300 83.700 1099.700 84.860 ;
        RECT 0.090 81.500 1099.700 83.700 ;
        RECT 0.090 80.340 0.700 81.500 ;
        RECT 4.300 80.340 1099.700 81.500 ;
        RECT 0.090 78.140 1099.700 80.340 ;
        RECT 0.090 76.980 1095.700 78.140 ;
        RECT 1099.300 76.980 1099.700 78.140 ;
        RECT 0.090 71.420 1099.700 76.980 ;
        RECT 0.090 70.260 0.700 71.420 ;
        RECT 4.300 70.260 1099.700 71.420 ;
        RECT 0.090 68.060 1099.700 70.260 ;
        RECT 0.090 66.900 1095.700 68.060 ;
        RECT 1099.300 66.900 1099.700 68.060 ;
        RECT 0.090 64.700 1099.700 66.900 ;
        RECT 0.090 63.540 0.700 64.700 ;
        RECT 4.300 63.540 1099.700 64.700 ;
        RECT 0.090 57.980 1099.700 63.540 ;
        RECT 0.090 56.820 1095.700 57.980 ;
        RECT 1099.300 56.820 1099.700 57.980 ;
        RECT 0.090 54.620 1099.700 56.820 ;
        RECT 0.090 53.460 0.700 54.620 ;
        RECT 4.300 53.460 1099.700 54.620 ;
        RECT 0.090 47.900 1099.700 53.460 ;
        RECT 0.090 46.740 1095.700 47.900 ;
        RECT 1099.300 46.740 1099.700 47.900 ;
        RECT 0.090 44.540 1099.700 46.740 ;
        RECT 0.090 43.380 0.700 44.540 ;
        RECT 4.300 43.380 1099.700 44.540 ;
        RECT 0.090 41.180 1099.700 43.380 ;
        RECT 0.090 40.020 1095.700 41.180 ;
        RECT 1099.300 40.020 1099.700 41.180 ;
        RECT 0.090 34.460 1099.700 40.020 ;
        RECT 0.090 33.300 0.700 34.460 ;
        RECT 4.300 33.300 1099.700 34.460 ;
        RECT 0.090 31.100 1099.700 33.300 ;
        RECT 0.090 29.940 1095.700 31.100 ;
        RECT 1099.300 29.940 1099.700 31.100 ;
        RECT 0.090 27.740 1099.700 29.940 ;
        RECT 0.090 26.580 0.700 27.740 ;
        RECT 4.300 26.580 1099.700 27.740 ;
        RECT 0.090 21.020 1099.700 26.580 ;
        RECT 0.090 19.860 1095.700 21.020 ;
        RECT 1099.300 19.860 1099.700 21.020 ;
        RECT 0.090 17.660 1099.700 19.860 ;
        RECT 0.090 16.500 0.700 17.660 ;
        RECT 4.300 16.500 1099.700 17.660 ;
        RECT 0.090 10.940 1099.700 16.500 ;
        RECT 0.090 9.780 1095.700 10.940 ;
        RECT 1099.300 9.780 1099.700 10.940 ;
        RECT 0.090 7.580 1099.700 9.780 ;
        RECT 0.090 6.420 0.700 7.580 ;
        RECT 4.300 6.420 1099.700 7.580 ;
        RECT 0.090 4.220 1099.700 6.420 ;
        RECT 0.090 3.500 1095.700 4.220 ;
        RECT 1099.300 3.500 1099.700 4.220 ;
  END
END tiny_user_project
END LIBRARY

