// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire net112;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net113;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net114;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net82;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net83;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net84;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net18;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net19;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net20;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net21;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net22;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net23;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net155;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net156;
 wire net184;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _004_ (.I(net3),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _005_ (.A1(net4),
    .A2(net14),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _006_ (.A1(net5),
    .A2(net13),
    .ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _007_ (.I(net7),
    .ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _008_ (.I(net11),
    .ZN(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _009_ (.I(net9),
    .ZN(net10));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _010_ (.A1(net6),
    .A2(net8),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _011_ (.A1(net6),
    .A2(net8),
    .B(net15),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _012_ (.A1(_002_),
    .A2(_003_),
    .ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _013_ (.A1(_000_),
    .A2(net2),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 _014_ (.D(net8),
    .RN(_000_),
    .SETN(_001_),
    .CLK(net1),
    .Q(net11));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _015_ (.D(net8),
    .CLK(net7),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_18 (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_19 (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_20 (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_21 (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[14]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[15]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[8]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[9]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output9 (.I(net9),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output10 (.I(net10),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output11 (.I(net11),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output12 (.I(net12),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output13 (.I(net13),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output14 (.I(net14),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output15 (.I(net15),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output16 (.I(net16),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_17 (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__014__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__013__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__004__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__006__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__011__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__010__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__015__CLK (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__007__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__015__D (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__014__D (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__011__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__010__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__009__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__008__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__006__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__005__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__011__B (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1936 ();
 assign io_oeb[0] = net111;
 assign io_oeb[10] = net121;
 assign io_oeb[11] = net122;
 assign io_oeb[12] = net123;
 assign io_oeb[13] = net124;
 assign io_oeb[14] = net125;
 assign io_oeb[15] = net126;
 assign io_oeb[16] = net127;
 assign io_oeb[17] = net128;
 assign io_oeb[18] = net129;
 assign io_oeb[19] = net130;
 assign io_oeb[1] = net112;
 assign io_oeb[20] = net131;
 assign io_oeb[21] = net132;
 assign io_oeb[22] = net133;
 assign io_oeb[23] = net134;
 assign io_oeb[24] = net135;
 assign io_oeb[25] = net136;
 assign io_oeb[26] = net137;
 assign io_oeb[27] = net138;
 assign io_oeb[28] = net139;
 assign io_oeb[29] = net140;
 assign io_oeb[2] = net113;
 assign io_oeb[30] = net141;
 assign io_oeb[31] = net142;
 assign io_oeb[32] = net143;
 assign io_oeb[33] = net144;
 assign io_oeb[34] = net145;
 assign io_oeb[35] = net146;
 assign io_oeb[36] = net147;
 assign io_oeb[37] = net148;
 assign io_oeb[3] = net114;
 assign io_oeb[4] = net115;
 assign io_oeb[5] = net116;
 assign io_oeb[6] = net117;
 assign io_oeb[7] = net118;
 assign io_oeb[8] = net119;
 assign io_oeb[9] = net120;
 assign io_out[0] = net81;
 assign io_out[10] = net91;
 assign io_out[11] = net92;
 assign io_out[12] = net93;
 assign io_out[13] = net94;
 assign io_out[14] = net95;
 assign io_out[15] = net96;
 assign io_out[1] = net82;
 assign io_out[24] = net97;
 assign io_out[25] = net98;
 assign io_out[26] = net99;
 assign io_out[27] = net100;
 assign io_out[28] = net101;
 assign io_out[29] = net102;
 assign io_out[2] = net83;
 assign io_out[30] = net103;
 assign io_out[31] = net104;
 assign io_out[32] = net105;
 assign io_out[33] = net106;
 assign io_out[34] = net107;
 assign io_out[35] = net108;
 assign io_out[36] = net109;
 assign io_out[37] = net110;
 assign io_out[3] = net84;
 assign io_out[4] = net85;
 assign io_out[5] = net86;
 assign io_out[6] = net87;
 assign io_out[7] = net88;
 assign io_out[8] = net89;
 assign io_out[9] = net90;
 assign la_data_out[0] = net17;
 assign la_data_out[10] = net27;
 assign la_data_out[11] = net28;
 assign la_data_out[12] = net29;
 assign la_data_out[13] = net30;
 assign la_data_out[14] = net31;
 assign la_data_out[15] = net32;
 assign la_data_out[16] = net33;
 assign la_data_out[17] = net34;
 assign la_data_out[18] = net35;
 assign la_data_out[19] = net36;
 assign la_data_out[1] = net18;
 assign la_data_out[20] = net37;
 assign la_data_out[21] = net38;
 assign la_data_out[22] = net39;
 assign la_data_out[23] = net40;
 assign la_data_out[24] = net41;
 assign la_data_out[25] = net42;
 assign la_data_out[26] = net43;
 assign la_data_out[27] = net44;
 assign la_data_out[28] = net45;
 assign la_data_out[29] = net46;
 assign la_data_out[2] = net19;
 assign la_data_out[30] = net47;
 assign la_data_out[31] = net48;
 assign la_data_out[32] = net49;
 assign la_data_out[33] = net50;
 assign la_data_out[34] = net51;
 assign la_data_out[35] = net52;
 assign la_data_out[36] = net53;
 assign la_data_out[37] = net54;
 assign la_data_out[38] = net55;
 assign la_data_out[39] = net56;
 assign la_data_out[3] = net20;
 assign la_data_out[40] = net57;
 assign la_data_out[41] = net58;
 assign la_data_out[42] = net59;
 assign la_data_out[43] = net60;
 assign la_data_out[44] = net61;
 assign la_data_out[45] = net62;
 assign la_data_out[46] = net63;
 assign la_data_out[47] = net64;
 assign la_data_out[48] = net65;
 assign la_data_out[49] = net66;
 assign la_data_out[4] = net21;
 assign la_data_out[50] = net67;
 assign la_data_out[51] = net68;
 assign la_data_out[52] = net69;
 assign la_data_out[53] = net70;
 assign la_data_out[54] = net71;
 assign la_data_out[55] = net72;
 assign la_data_out[56] = net73;
 assign la_data_out[57] = net74;
 assign la_data_out[58] = net75;
 assign la_data_out[59] = net76;
 assign la_data_out[5] = net22;
 assign la_data_out[60] = net77;
 assign la_data_out[61] = net78;
 assign la_data_out[62] = net79;
 assign la_data_out[63] = net80;
 assign la_data_out[6] = net23;
 assign la_data_out[7] = net24;
 assign la_data_out[8] = net25;
 assign la_data_out[9] = net26;
 assign user_irq[0] = net149;
 assign user_irq[1] = net150;
 assign user_irq[2] = net151;
 assign wbs_ack_o = net152;
 assign wbs_dat_o[0] = net153;
 assign wbs_dat_o[10] = net163;
 assign wbs_dat_o[11] = net164;
 assign wbs_dat_o[12] = net165;
 assign wbs_dat_o[13] = net166;
 assign wbs_dat_o[14] = net167;
 assign wbs_dat_o[15] = net168;
 assign wbs_dat_o[16] = net169;
 assign wbs_dat_o[17] = net170;
 assign wbs_dat_o[18] = net171;
 assign wbs_dat_o[19] = net172;
 assign wbs_dat_o[1] = net154;
 assign wbs_dat_o[20] = net173;
 assign wbs_dat_o[21] = net174;
 assign wbs_dat_o[22] = net175;
 assign wbs_dat_o[23] = net176;
 assign wbs_dat_o[24] = net177;
 assign wbs_dat_o[25] = net178;
 assign wbs_dat_o[26] = net179;
 assign wbs_dat_o[27] = net180;
 assign wbs_dat_o[28] = net181;
 assign wbs_dat_o[29] = net182;
 assign wbs_dat_o[2] = net155;
 assign wbs_dat_o[30] = net183;
 assign wbs_dat_o[31] = net184;
 assign wbs_dat_o[3] = net156;
 assign wbs_dat_o[4] = net157;
 assign wbs_dat_o[5] = net158;
 assign wbs_dat_o[6] = net159;
 assign wbs_dat_o[7] = net160;
 assign wbs_dat_o[8] = net161;
 assign wbs_dat_o[9] = net162;
endmodule

