VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 3000.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 33.320 3004.800 34.440 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2032.520 3004.800 2033.640 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2232.440 3004.800 2233.560 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2432.360 3004.800 2433.480 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2632.280 3004.800 2633.400 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2832.200 3004.800 2833.320 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2940.840 2997.600 2941.960 3004.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2608.200 2997.600 2609.320 3004.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2275.560 2997.600 2276.680 3004.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1942.920 2997.600 1944.040 3004.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1610.280 2997.600 1611.400 3004.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 233.240 3004.800 234.360 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1277.640 2997.600 1278.760 3004.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 945.000 2997.600 946.120 3004.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 612.360 2997.600 613.480 3004.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.720 2997.600 280.840 3004.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2957.080 2.400 2958.200 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2743.720 2.400 2744.840 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2530.360 2.400 2531.480 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2317.000 2.400 2318.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2103.640 2.400 2104.760 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1890.280 2.400 1891.400 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 433.160 3004.800 434.280 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1676.920 2.400 1678.040 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1463.560 2.400 1464.680 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1250.200 2.400 1251.320 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1036.840 2.400 1037.960 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 823.480 2.400 824.600 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 610.120 2.400 611.240 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 396.760 2.400 397.880 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 183.400 2.400 184.520 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 633.080 3004.800 634.200 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 833.000 3004.800 834.120 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1032.920 3004.800 1034.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1232.840 3004.800 1233.960 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1432.760 3004.800 1433.880 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1632.680 3004.800 1633.800 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1832.600 3004.800 1833.720 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 166.600 3004.800 167.720 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2165.800 3004.800 2166.920 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2365.720 3004.800 2366.840 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2565.640 3004.800 2566.760 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2765.560 3004.800 2766.680 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2965.480 3004.800 2966.600 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2719.080 2997.600 2720.200 3004.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2386.440 2997.600 2387.560 3004.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2053.800 2997.600 2054.920 3004.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1721.160 2997.600 1722.280 3004.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1388.520 2997.600 1389.640 3004.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 366.520 3004.800 367.640 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1055.880 2997.600 1057.000 3004.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 723.240 2997.600 724.360 3004.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.600 2997.600 391.720 3004.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.960 2997.600 59.080 3004.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2814.840 2.400 2815.960 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2601.480 2.400 2602.600 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2388.120 2.400 2389.240 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2174.760 2.400 2175.880 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1961.400 2.400 1962.520 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1748.040 2.400 1749.160 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 566.440 3004.800 567.560 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1534.680 2.400 1535.800 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1321.320 2.400 1322.440 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1107.960 2.400 1109.080 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 894.600 2.400 895.720 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 681.240 2.400 682.360 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 467.880 2.400 469.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 254.520 2.400 255.640 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 41.160 2.400 42.280 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 766.360 3004.800 767.480 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 966.280 3004.800 967.400 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1166.200 3004.800 1167.320 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1366.120 3004.800 1367.240 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1566.040 3004.800 1567.160 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1765.960 3004.800 1767.080 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1965.880 3004.800 1967.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 99.960 3004.800 101.080 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2099.160 3004.800 2100.280 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2299.080 3004.800 2300.200 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2499.000 3004.800 2500.120 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2698.920 3004.800 2700.040 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 2898.840 3004.800 2899.960 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2829.960 2997.600 2831.080 3004.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2497.320 2997.600 2498.440 3004.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2164.680 2997.600 2165.800 3004.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1832.040 2997.600 1833.160 3004.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1499.400 2997.600 1500.520 3004.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 299.880 3004.800 301.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1166.760 2997.600 1167.880 3004.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 834.120 2997.600 835.240 3004.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 501.480 2997.600 502.600 3004.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.840 2997.600 169.960 3004.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2885.960 2.400 2887.080 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2672.600 2.400 2673.720 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2459.240 2.400 2460.360 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2245.880 2.400 2247.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 2032.520 2.400 2033.640 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1819.160 2.400 1820.280 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 499.800 3004.800 500.920 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1605.800 2.400 1606.920 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1392.440 2.400 1393.560 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 1179.080 2.400 1180.200 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 965.720 2.400 966.840 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 752.360 2.400 753.480 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 539.000 2.400 540.120 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 325.640 2.400 326.760 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.800 112.280 2.400 113.400 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 699.720 3004.800 700.840 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 899.640 3004.800 900.760 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1099.560 3004.800 1100.680 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1299.480 3004.800 1300.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1499.400 3004.800 1500.520 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1699.320 3004.800 1700.440 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2997.600 1899.240 3004.800 1900.360 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1075.480 -4.800 1076.600 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1361.080 -4.800 1362.200 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1389.640 -4.800 1390.760 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1418.200 -4.800 1419.320 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1446.760 -4.800 1447.880 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1475.320 -4.800 1476.440 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1503.880 -4.800 1505.000 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1532.440 -4.800 1533.560 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1561.000 -4.800 1562.120 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1589.560 -4.800 1590.680 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1618.120 -4.800 1619.240 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1104.040 -4.800 1105.160 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1646.680 -4.800 1647.800 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1675.240 -4.800 1676.360 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1703.800 -4.800 1704.920 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1732.360 -4.800 1733.480 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1760.920 -4.800 1762.040 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1789.480 -4.800 1790.600 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1818.040 -4.800 1819.160 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1846.600 -4.800 1847.720 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1875.160 -4.800 1876.280 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1903.720 -4.800 1904.840 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1132.600 -4.800 1133.720 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1932.280 -4.800 1933.400 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1960.840 -4.800 1961.960 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1989.400 -4.800 1990.520 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2017.960 -4.800 2019.080 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2046.520 -4.800 2047.640 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2075.080 -4.800 2076.200 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2103.640 -4.800 2104.760 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2132.200 -4.800 2133.320 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2160.760 -4.800 2161.880 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2189.320 -4.800 2190.440 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1161.160 -4.800 1162.280 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2217.880 -4.800 2219.000 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2246.440 -4.800 2247.560 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2275.000 -4.800 2276.120 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2303.560 -4.800 2304.680 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2332.120 -4.800 2333.240 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2360.680 -4.800 2361.800 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2389.240 -4.800 2390.360 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2417.800 -4.800 2418.920 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2446.360 -4.800 2447.480 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2474.920 -4.800 2476.040 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1189.720 -4.800 1190.840 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2503.480 -4.800 2504.600 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2532.040 -4.800 2533.160 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2560.600 -4.800 2561.720 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2589.160 -4.800 2590.280 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2617.720 -4.800 2618.840 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2646.280 -4.800 2647.400 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2674.840 -4.800 2675.960 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2703.400 -4.800 2704.520 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2731.960 -4.800 2733.080 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2760.520 -4.800 2761.640 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1218.280 -4.800 1219.400 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2789.080 -4.800 2790.200 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2817.640 -4.800 2818.760 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2846.200 -4.800 2847.320 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2874.760 -4.800 2875.880 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1246.840 -4.800 1247.960 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1275.400 -4.800 1276.520 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1303.960 -4.800 1305.080 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1332.520 -4.800 1333.640 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1085.000 -4.800 1086.120 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1370.600 -4.800 1371.720 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1399.160 -4.800 1400.280 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1427.720 -4.800 1428.840 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1456.280 -4.800 1457.400 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1484.840 -4.800 1485.960 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1513.400 -4.800 1514.520 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1541.960 -4.800 1543.080 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1570.520 -4.800 1571.640 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1599.080 -4.800 1600.200 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1627.640 -4.800 1628.760 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1113.560 -4.800 1114.680 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1656.200 -4.800 1657.320 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1684.760 -4.800 1685.880 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1713.320 -4.800 1714.440 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1741.880 -4.800 1743.000 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1770.440 -4.800 1771.560 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1799.000 -4.800 1800.120 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1827.560 -4.800 1828.680 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1856.120 -4.800 1857.240 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1884.680 -4.800 1885.800 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1913.240 -4.800 1914.360 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1142.120 -4.800 1143.240 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1941.800 -4.800 1942.920 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1970.360 -4.800 1971.480 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1998.920 -4.800 2000.040 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2027.480 -4.800 2028.600 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2056.040 -4.800 2057.160 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2084.600 -4.800 2085.720 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2113.160 -4.800 2114.280 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2141.720 -4.800 2142.840 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2170.280 -4.800 2171.400 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2198.840 -4.800 2199.960 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1170.680 -4.800 1171.800 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2227.400 -4.800 2228.520 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2255.960 -4.800 2257.080 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2284.520 -4.800 2285.640 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2313.080 -4.800 2314.200 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2341.640 -4.800 2342.760 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2370.200 -4.800 2371.320 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2398.760 -4.800 2399.880 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2427.320 -4.800 2428.440 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2455.880 -4.800 2457.000 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2484.440 -4.800 2485.560 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1199.240 -4.800 1200.360 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2513.000 -4.800 2514.120 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2541.560 -4.800 2542.680 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2570.120 -4.800 2571.240 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2598.680 -4.800 2599.800 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2627.240 -4.800 2628.360 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2655.800 -4.800 2656.920 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2684.360 -4.800 2685.480 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2712.920 -4.800 2714.040 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2741.480 -4.800 2742.600 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2770.040 -4.800 2771.160 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1227.800 -4.800 1228.920 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2798.600 -4.800 2799.720 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2827.160 -4.800 2828.280 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2855.720 -4.800 2856.840 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2884.280 -4.800 2885.400 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1256.360 -4.800 1257.480 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1284.920 -4.800 1286.040 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1313.480 -4.800 1314.600 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1342.040 -4.800 1343.160 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1094.520 -4.800 1095.640 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1380.120 -4.800 1381.240 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1408.680 -4.800 1409.800 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1437.240 -4.800 1438.360 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1465.800 -4.800 1466.920 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1494.360 -4.800 1495.480 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1522.920 -4.800 1524.040 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1551.480 -4.800 1552.600 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1580.040 -4.800 1581.160 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1608.600 -4.800 1609.720 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1637.160 -4.800 1638.280 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1123.080 -4.800 1124.200 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1665.720 -4.800 1666.840 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1694.280 -4.800 1695.400 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1722.840 -4.800 1723.960 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1751.400 -4.800 1752.520 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1779.960 -4.800 1781.080 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1808.520 -4.800 1809.640 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1837.080 -4.800 1838.200 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1865.640 -4.800 1866.760 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1894.200 -4.800 1895.320 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1922.760 -4.800 1923.880 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1151.640 -4.800 1152.760 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1951.320 -4.800 1952.440 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1979.880 -4.800 1981.000 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2008.440 -4.800 2009.560 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2037.000 -4.800 2038.120 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2065.560 -4.800 2066.680 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2094.120 -4.800 2095.240 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2122.680 -4.800 2123.800 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2151.240 -4.800 2152.360 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2179.800 -4.800 2180.920 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2208.360 -4.800 2209.480 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1180.200 -4.800 1181.320 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2236.920 -4.800 2238.040 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2265.480 -4.800 2266.600 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2294.040 -4.800 2295.160 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2322.600 -4.800 2323.720 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2351.160 -4.800 2352.280 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2379.720 -4.800 2380.840 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2408.280 -4.800 2409.400 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2436.840 -4.800 2437.960 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2465.400 -4.800 2466.520 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2493.960 -4.800 2495.080 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1208.760 -4.800 1209.880 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2522.520 -4.800 2523.640 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2551.080 -4.800 2552.200 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2579.640 -4.800 2580.760 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2608.200 -4.800 2609.320 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2636.760 -4.800 2637.880 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2665.320 -4.800 2666.440 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2693.880 -4.800 2695.000 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2722.440 -4.800 2723.560 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2751.000 -4.800 2752.120 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2779.560 -4.800 2780.680 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1237.320 -4.800 1238.440 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2808.120 -4.800 2809.240 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2836.680 -4.800 2837.800 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2865.240 -4.800 2866.360 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2893.800 -4.800 2894.920 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1265.880 -4.800 1267.000 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1294.440 -4.800 1295.560 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1323.000 -4.800 1324.120 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1351.560 -4.800 1352.680 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2903.320 -4.800 2904.440 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2912.840 -4.800 2913.960 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2922.360 -4.800 2923.480 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2931.880 -4.800 2933.000 2.400 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 4.740 6.420 7.840 2992.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.740 6.420 2995.180 9.520 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.740 2989.280 2995.180 2992.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2992.080 6.420 2995.180 2992.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 25.290 1.620 28.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 115.290 1.620 118.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 205.290 1.620 208.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 295.290 1.620 298.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 385.290 1.620 388.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 475.290 1.620 478.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 565.290 1.620 568.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 655.290 1.620 658.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 745.290 1.620 748.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 835.290 1.620 838.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 925.290 1.620 928.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1015.290 1.620 1018.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1105.290 1.620 1108.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1195.290 1.620 1198.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1285.290 1.620 1288.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1375.290 1.620 1378.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1465.290 1.620 1468.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1555.290 1.620 1558.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1645.290 1.620 1648.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1735.290 1.620 1738.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1825.290 1.620 1828.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1915.290 1.620 1918.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2005.290 1.620 2008.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.290 1.620 2098.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2185.290 1.620 2188.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2275.290 1.620 2278.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2365.290 1.620 2368.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2455.290 1.620 2458.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2545.290 1.620 2548.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2635.290 1.620 2638.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2725.290 1.620 2728.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2815.290 1.620 2818.390 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2905.290 1.620 2908.390 2997.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 26.970 2999.980 30.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 116.970 2999.980 120.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 206.970 2999.980 210.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 296.970 2999.980 300.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 386.970 2999.980 390.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 476.970 2999.980 480.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 566.970 2999.980 570.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 656.970 2999.980 660.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 746.970 2999.980 750.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 836.970 2999.980 840.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 926.970 2999.980 930.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1016.970 2999.980 1020.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1106.970 2999.980 1110.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1196.970 2999.980 1200.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1286.970 2999.980 1290.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1376.970 2999.980 1380.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1466.970 2999.980 1470.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1556.970 2999.980 1560.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1646.970 2999.980 1650.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1736.970 2999.980 1740.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1826.970 2999.980 1830.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1916.970 2999.980 1920.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2006.970 2999.980 2010.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2096.970 2999.980 2100.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2186.970 2999.980 2190.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2276.970 2999.980 2280.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2366.970 2999.980 2370.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2456.970 2999.980 2460.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2546.970 2999.980 2550.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2636.970 2999.980 2640.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2726.970 2999.980 2730.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2816.970 2999.980 2820.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2906.970 2999.980 2910.070 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -0.060 1.620 3.040 2997.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1.620 2999.980 4.720 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2994.080 2999.980 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2996.880 1.620 2999.980 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.890 1.620 46.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 133.890 1.620 136.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 223.890 1.620 226.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 313.890 1.620 316.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 403.890 1.620 406.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 493.890 1.620 496.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 583.890 1.620 586.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 673.890 1.620 676.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 763.890 1.620 766.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 853.890 1.620 856.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.890 1.620 946.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1033.890 1.620 1036.990 555.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1033.890 1344.580 1036.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1123.890 1.620 1126.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1213.890 1.620 1216.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1303.890 1.620 1306.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1393.890 1.620 1396.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1483.890 1.620 1486.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1573.890 1.620 1576.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1663.890 1.620 1666.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1753.890 1.620 1756.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1843.890 1.620 1846.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1933.890 1.620 1936.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2023.890 1.620 2026.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2113.890 1.620 2116.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2203.890 1.620 2206.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2293.890 1.620 2296.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2383.890 1.620 2386.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2473.890 1.620 2476.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2563.890 1.620 2566.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2653.890 1.620 2656.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2743.890 1.620 2746.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2833.890 1.620 2836.990 2997.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2923.890 1.620 2926.990 2997.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 56.970 2999.980 60.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 146.970 2999.980 150.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 236.970 2999.980 240.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 326.970 2999.980 330.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 416.970 2999.980 420.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 506.970 2999.980 510.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 596.970 2999.980 600.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 686.970 2999.980 690.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 776.970 2999.980 780.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 866.970 2999.980 870.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 956.970 2999.980 960.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1046.970 2999.980 1050.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1136.970 2999.980 1140.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1226.970 2999.980 1230.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1316.970 2999.980 1320.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1406.970 2999.980 1410.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1496.970 2999.980 1500.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1586.970 2999.980 1590.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1676.970 2999.980 1680.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1766.970 2999.980 1770.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1856.970 2999.980 1860.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 1946.970 2999.980 1950.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2036.970 2999.980 2040.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2126.970 2999.980 2130.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2216.970 2999.980 2220.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2306.970 2999.980 2310.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2396.970 2999.980 2400.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2486.970 2999.980 2490.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2576.970 2999.980 2580.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2666.970 2999.980 2670.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2756.970 2999.980 2760.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2846.970 2999.980 2850.070 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.060 2936.970 2999.980 2940.070 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.360 -4.800 67.480 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 75.880 -4.800 77.000 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 85.400 -4.800 86.520 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.480 -4.800 124.600 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 447.160 -4.800 448.280 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 475.720 -4.800 476.840 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.280 -4.800 505.400 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.840 -4.800 533.960 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.400 -4.800 562.520 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 589.960 -4.800 591.080 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.520 -4.800 619.640 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 647.080 -4.800 648.200 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.640 -4.800 676.760 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 704.200 -4.800 705.320 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.560 -4.800 162.680 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.760 -4.800 733.880 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 761.320 -4.800 762.440 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.880 -4.800 791.000 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 818.440 -4.800 819.560 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 847.000 -4.800 848.120 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 875.560 -4.800 876.680 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 904.120 -4.800 905.240 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 932.680 -4.800 933.800 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 961.240 -4.800 962.360 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 989.800 -4.800 990.920 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.640 -4.800 200.760 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1018.360 -4.800 1019.480 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1046.920 -4.800 1048.040 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 237.720 -4.800 238.840 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.800 -4.800 276.920 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.360 -4.800 305.480 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.920 -4.800 334.040 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 361.480 -4.800 362.600 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.040 -4.800 391.160 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.600 -4.800 419.720 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.920 -4.800 96.040 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.000 -4.800 134.120 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.680 -4.800 457.800 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 485.240 -4.800 486.360 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 513.800 -4.800 514.920 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.360 -4.800 543.480 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 570.920 -4.800 572.040 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.480 -4.800 600.600 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.040 -4.800 629.160 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 656.600 -4.800 657.720 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.160 -4.800 686.280 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 713.720 -4.800 714.840 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.080 -4.800 172.200 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.280 -4.800 743.400 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 770.840 -4.800 771.960 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.400 -4.800 800.520 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 827.960 -4.800 829.080 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.520 -4.800 857.640 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 885.080 -4.800 886.200 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 913.640 -4.800 914.760 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 942.200 -4.800 943.320 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 970.760 -4.800 971.880 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 999.320 -4.800 1000.440 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.160 -4.800 210.280 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1027.880 -4.800 1029.000 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1056.440 -4.800 1057.560 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.240 -4.800 248.360 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.320 -4.800 286.440 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.880 -4.800 315.000 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.440 -4.800 343.560 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.000 -4.800 372.120 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.560 -4.800 400.680 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 428.120 -4.800 429.240 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.520 -4.800 143.640 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 466.200 -4.800 467.320 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 494.760 -4.800 495.880 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.320 -4.800 524.440 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.880 -4.800 553.000 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 580.440 -4.800 581.560 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 609.000 -4.800 610.120 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 637.560 -4.800 638.680 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 666.120 -4.800 667.240 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 694.680 -4.800 695.800 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 723.240 -4.800 724.360 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.600 -4.800 181.720 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 751.800 -4.800 752.920 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 780.360 -4.800 781.480 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 808.920 -4.800 810.040 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 837.480 -4.800 838.600 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 866.040 -4.800 867.160 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 894.600 -4.800 895.720 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 923.160 -4.800 924.280 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 951.720 -4.800 952.840 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 980.280 -4.800 981.400 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1008.840 -4.800 1009.960 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.680 -4.800 219.800 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1037.400 -4.800 1038.520 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1065.960 -4.800 1067.080 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.760 -4.800 257.880 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.840 -4.800 295.960 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.400 -4.800 324.520 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.960 -4.800 353.080 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.520 -4.800 381.640 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.080 -4.800 410.200 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.640 -4.800 438.760 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 152.040 -4.800 153.160 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.120 -4.800 191.240 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.200 -4.800 229.320 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.280 -4.800 267.400 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.440 -4.800 105.560 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 -4.800 115.080 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 406.720 527.670 1493.120 1334.970 ;
      LAYER Metal2 ;
        RECT 12.460 2997.300 57.660 2998.100 ;
        RECT 59.380 2997.300 168.540 2998.100 ;
        RECT 170.260 2997.300 279.420 2998.100 ;
        RECT 281.140 2997.300 390.300 2998.100 ;
        RECT 392.020 2997.300 501.180 2998.100 ;
        RECT 502.900 2997.300 612.060 2998.100 ;
        RECT 613.780 2997.300 722.940 2998.100 ;
        RECT 724.660 2997.300 833.820 2998.100 ;
        RECT 835.540 2997.300 944.700 2998.100 ;
        RECT 946.420 2997.300 1055.580 2998.100 ;
        RECT 1057.300 2997.300 1166.460 2998.100 ;
        RECT 1168.180 2997.300 1277.340 2998.100 ;
        RECT 1279.060 2997.300 1388.220 2998.100 ;
        RECT 1389.940 2997.300 1499.100 2998.100 ;
        RECT 1500.820 2997.300 1609.980 2998.100 ;
        RECT 1611.700 2997.300 1720.860 2998.100 ;
        RECT 1722.580 2997.300 1831.740 2998.100 ;
        RECT 1833.460 2997.300 1942.620 2998.100 ;
        RECT 1944.340 2997.300 2053.500 2998.100 ;
        RECT 2055.220 2997.300 2164.380 2998.100 ;
        RECT 2166.100 2997.300 2275.260 2998.100 ;
        RECT 2276.980 2997.300 2386.140 2998.100 ;
        RECT 2387.860 2997.300 2497.020 2998.100 ;
        RECT 2498.740 2997.300 2607.900 2998.100 ;
        RECT 2609.620 2997.300 2718.780 2998.100 ;
        RECT 2720.500 2997.300 2829.660 2998.100 ;
        RECT 2831.380 2997.300 2940.540 2998.100 ;
        RECT 2942.260 2997.300 2992.500 2998.100 ;
        RECT 12.460 2.700 2992.500 2997.300 ;
        RECT 12.460 0.090 66.060 2.700 ;
        RECT 67.780 0.090 75.580 2.700 ;
        RECT 77.300 0.090 85.100 2.700 ;
        RECT 86.820 0.090 94.620 2.700 ;
        RECT 96.340 0.090 104.140 2.700 ;
        RECT 105.860 0.090 113.660 2.700 ;
        RECT 115.380 0.090 123.180 2.700 ;
        RECT 124.900 0.090 132.700 2.700 ;
        RECT 134.420 0.090 142.220 2.700 ;
        RECT 143.940 0.090 151.740 2.700 ;
        RECT 153.460 0.090 161.260 2.700 ;
        RECT 162.980 0.090 170.780 2.700 ;
        RECT 172.500 0.090 180.300 2.700 ;
        RECT 182.020 0.090 189.820 2.700 ;
        RECT 191.540 0.090 199.340 2.700 ;
        RECT 201.060 0.090 208.860 2.700 ;
        RECT 210.580 0.090 218.380 2.700 ;
        RECT 220.100 0.090 227.900 2.700 ;
        RECT 229.620 0.090 237.420 2.700 ;
        RECT 239.140 0.090 246.940 2.700 ;
        RECT 248.660 0.090 256.460 2.700 ;
        RECT 258.180 0.090 265.980 2.700 ;
        RECT 267.700 0.090 275.500 2.700 ;
        RECT 277.220 0.090 285.020 2.700 ;
        RECT 286.740 0.090 294.540 2.700 ;
        RECT 296.260 0.090 304.060 2.700 ;
        RECT 305.780 0.090 313.580 2.700 ;
        RECT 315.300 0.090 323.100 2.700 ;
        RECT 324.820 0.090 332.620 2.700 ;
        RECT 334.340 0.090 342.140 2.700 ;
        RECT 343.860 0.090 351.660 2.700 ;
        RECT 353.380 0.090 361.180 2.700 ;
        RECT 362.900 0.090 370.700 2.700 ;
        RECT 372.420 0.090 380.220 2.700 ;
        RECT 381.940 0.090 389.740 2.700 ;
        RECT 391.460 0.090 399.260 2.700 ;
        RECT 400.980 0.090 408.780 2.700 ;
        RECT 410.500 0.090 418.300 2.700 ;
        RECT 420.020 0.090 427.820 2.700 ;
        RECT 429.540 0.090 437.340 2.700 ;
        RECT 439.060 0.090 446.860 2.700 ;
        RECT 448.580 0.090 456.380 2.700 ;
        RECT 458.100 0.090 465.900 2.700 ;
        RECT 467.620 0.090 475.420 2.700 ;
        RECT 477.140 0.090 484.940 2.700 ;
        RECT 486.660 0.090 494.460 2.700 ;
        RECT 496.180 0.090 503.980 2.700 ;
        RECT 505.700 0.090 513.500 2.700 ;
        RECT 515.220 0.090 523.020 2.700 ;
        RECT 524.740 0.090 532.540 2.700 ;
        RECT 534.260 0.090 542.060 2.700 ;
        RECT 543.780 0.090 551.580 2.700 ;
        RECT 553.300 0.090 561.100 2.700 ;
        RECT 562.820 0.090 570.620 2.700 ;
        RECT 572.340 0.090 580.140 2.700 ;
        RECT 581.860 0.090 589.660 2.700 ;
        RECT 591.380 0.090 599.180 2.700 ;
        RECT 600.900 0.090 608.700 2.700 ;
        RECT 610.420 0.090 618.220 2.700 ;
        RECT 619.940 0.090 627.740 2.700 ;
        RECT 629.460 0.090 637.260 2.700 ;
        RECT 638.980 0.090 646.780 2.700 ;
        RECT 648.500 0.090 656.300 2.700 ;
        RECT 658.020 0.090 665.820 2.700 ;
        RECT 667.540 0.090 675.340 2.700 ;
        RECT 677.060 0.090 684.860 2.700 ;
        RECT 686.580 0.090 694.380 2.700 ;
        RECT 696.100 0.090 703.900 2.700 ;
        RECT 705.620 0.090 713.420 2.700 ;
        RECT 715.140 0.090 722.940 2.700 ;
        RECT 724.660 0.090 732.460 2.700 ;
        RECT 734.180 0.090 741.980 2.700 ;
        RECT 743.700 0.090 751.500 2.700 ;
        RECT 753.220 0.090 761.020 2.700 ;
        RECT 762.740 0.090 770.540 2.700 ;
        RECT 772.260 0.090 780.060 2.700 ;
        RECT 781.780 0.090 789.580 2.700 ;
        RECT 791.300 0.090 799.100 2.700 ;
        RECT 800.820 0.090 808.620 2.700 ;
        RECT 810.340 0.090 818.140 2.700 ;
        RECT 819.860 0.090 827.660 2.700 ;
        RECT 829.380 0.090 837.180 2.700 ;
        RECT 838.900 0.090 846.700 2.700 ;
        RECT 848.420 0.090 856.220 2.700 ;
        RECT 857.940 0.090 865.740 2.700 ;
        RECT 867.460 0.090 875.260 2.700 ;
        RECT 876.980 0.090 884.780 2.700 ;
        RECT 886.500 0.090 894.300 2.700 ;
        RECT 896.020 0.090 903.820 2.700 ;
        RECT 905.540 0.090 913.340 2.700 ;
        RECT 915.060 0.090 922.860 2.700 ;
        RECT 924.580 0.090 932.380 2.700 ;
        RECT 934.100 0.090 941.900 2.700 ;
        RECT 943.620 0.090 951.420 2.700 ;
        RECT 953.140 0.090 960.940 2.700 ;
        RECT 962.660 0.090 970.460 2.700 ;
        RECT 972.180 0.090 979.980 2.700 ;
        RECT 981.700 0.090 989.500 2.700 ;
        RECT 991.220 0.090 999.020 2.700 ;
        RECT 1000.740 0.090 1008.540 2.700 ;
        RECT 1010.260 0.090 1018.060 2.700 ;
        RECT 1019.780 0.090 1027.580 2.700 ;
        RECT 1029.300 0.090 1037.100 2.700 ;
        RECT 1038.820 0.090 1046.620 2.700 ;
        RECT 1048.340 0.090 1056.140 2.700 ;
        RECT 1057.860 0.090 1065.660 2.700 ;
        RECT 1067.380 0.090 1075.180 2.700 ;
        RECT 1076.900 0.090 1084.700 2.700 ;
        RECT 1086.420 0.090 1094.220 2.700 ;
        RECT 1095.940 0.090 1103.740 2.700 ;
        RECT 1105.460 0.090 1113.260 2.700 ;
        RECT 1114.980 0.090 1122.780 2.700 ;
        RECT 1124.500 0.090 1132.300 2.700 ;
        RECT 1134.020 0.090 1141.820 2.700 ;
        RECT 1143.540 0.090 1151.340 2.700 ;
        RECT 1153.060 0.090 1160.860 2.700 ;
        RECT 1162.580 0.090 1170.380 2.700 ;
        RECT 1172.100 0.090 1179.900 2.700 ;
        RECT 1181.620 0.090 1189.420 2.700 ;
        RECT 1191.140 0.090 1198.940 2.700 ;
        RECT 1200.660 0.090 1208.460 2.700 ;
        RECT 1210.180 0.090 1217.980 2.700 ;
        RECT 1219.700 0.090 1227.500 2.700 ;
        RECT 1229.220 0.090 1237.020 2.700 ;
        RECT 1238.740 0.090 1246.540 2.700 ;
        RECT 1248.260 0.090 1256.060 2.700 ;
        RECT 1257.780 0.090 1265.580 2.700 ;
        RECT 1267.300 0.090 1275.100 2.700 ;
        RECT 1276.820 0.090 1284.620 2.700 ;
        RECT 1286.340 0.090 1294.140 2.700 ;
        RECT 1295.860 0.090 1303.660 2.700 ;
        RECT 1305.380 0.090 1313.180 2.700 ;
        RECT 1314.900 0.090 1322.700 2.700 ;
        RECT 1324.420 0.090 1332.220 2.700 ;
        RECT 1333.940 0.090 1341.740 2.700 ;
        RECT 1343.460 0.090 1351.260 2.700 ;
        RECT 1352.980 0.090 1360.780 2.700 ;
        RECT 1362.500 0.090 1370.300 2.700 ;
        RECT 1372.020 0.090 1379.820 2.700 ;
        RECT 1381.540 0.090 1389.340 2.700 ;
        RECT 1391.060 0.090 1398.860 2.700 ;
        RECT 1400.580 0.090 1408.380 2.700 ;
        RECT 1410.100 0.090 1417.900 2.700 ;
        RECT 1419.620 0.090 1427.420 2.700 ;
        RECT 1429.140 0.090 1436.940 2.700 ;
        RECT 1438.660 0.090 1446.460 2.700 ;
        RECT 1448.180 0.090 1455.980 2.700 ;
        RECT 1457.700 0.090 1465.500 2.700 ;
        RECT 1467.220 0.090 1475.020 2.700 ;
        RECT 1476.740 0.090 1484.540 2.700 ;
        RECT 1486.260 0.090 1494.060 2.700 ;
        RECT 1495.780 0.090 1503.580 2.700 ;
        RECT 1505.300 0.090 1513.100 2.700 ;
        RECT 1514.820 0.090 1522.620 2.700 ;
        RECT 1524.340 0.090 1532.140 2.700 ;
        RECT 1533.860 0.090 1541.660 2.700 ;
        RECT 1543.380 0.090 1551.180 2.700 ;
        RECT 1552.900 0.090 1560.700 2.700 ;
        RECT 1562.420 0.090 1570.220 2.700 ;
        RECT 1571.940 0.090 1579.740 2.700 ;
        RECT 1581.460 0.090 1589.260 2.700 ;
        RECT 1590.980 0.090 1598.780 2.700 ;
        RECT 1600.500 0.090 1608.300 2.700 ;
        RECT 1610.020 0.090 1617.820 2.700 ;
        RECT 1619.540 0.090 1627.340 2.700 ;
        RECT 1629.060 0.090 1636.860 2.700 ;
        RECT 1638.580 0.090 1646.380 2.700 ;
        RECT 1648.100 0.090 1655.900 2.700 ;
        RECT 1657.620 0.090 1665.420 2.700 ;
        RECT 1667.140 0.090 1674.940 2.700 ;
        RECT 1676.660 0.090 1684.460 2.700 ;
        RECT 1686.180 0.090 1693.980 2.700 ;
        RECT 1695.700 0.090 1703.500 2.700 ;
        RECT 1705.220 0.090 1713.020 2.700 ;
        RECT 1714.740 0.090 1722.540 2.700 ;
        RECT 1724.260 0.090 1732.060 2.700 ;
        RECT 1733.780 0.090 1741.580 2.700 ;
        RECT 1743.300 0.090 1751.100 2.700 ;
        RECT 1752.820 0.090 1760.620 2.700 ;
        RECT 1762.340 0.090 1770.140 2.700 ;
        RECT 1771.860 0.090 1779.660 2.700 ;
        RECT 1781.380 0.090 1789.180 2.700 ;
        RECT 1790.900 0.090 1798.700 2.700 ;
        RECT 1800.420 0.090 1808.220 2.700 ;
        RECT 1809.940 0.090 1817.740 2.700 ;
        RECT 1819.460 0.090 1827.260 2.700 ;
        RECT 1828.980 0.090 1836.780 2.700 ;
        RECT 1838.500 0.090 1846.300 2.700 ;
        RECT 1848.020 0.090 1855.820 2.700 ;
        RECT 1857.540 0.090 1865.340 2.700 ;
        RECT 1867.060 0.090 1874.860 2.700 ;
        RECT 1876.580 0.090 1884.380 2.700 ;
        RECT 1886.100 0.090 1893.900 2.700 ;
        RECT 1895.620 0.090 1903.420 2.700 ;
        RECT 1905.140 0.090 1912.940 2.700 ;
        RECT 1914.660 0.090 1922.460 2.700 ;
        RECT 1924.180 0.090 1931.980 2.700 ;
        RECT 1933.700 0.090 1941.500 2.700 ;
        RECT 1943.220 0.090 1951.020 2.700 ;
        RECT 1952.740 0.090 1960.540 2.700 ;
        RECT 1962.260 0.090 1970.060 2.700 ;
        RECT 1971.780 0.090 1979.580 2.700 ;
        RECT 1981.300 0.090 1989.100 2.700 ;
        RECT 1990.820 0.090 1998.620 2.700 ;
        RECT 2000.340 0.090 2008.140 2.700 ;
        RECT 2009.860 0.090 2017.660 2.700 ;
        RECT 2019.380 0.090 2027.180 2.700 ;
        RECT 2028.900 0.090 2036.700 2.700 ;
        RECT 2038.420 0.090 2046.220 2.700 ;
        RECT 2047.940 0.090 2055.740 2.700 ;
        RECT 2057.460 0.090 2065.260 2.700 ;
        RECT 2066.980 0.090 2074.780 2.700 ;
        RECT 2076.500 0.090 2084.300 2.700 ;
        RECT 2086.020 0.090 2093.820 2.700 ;
        RECT 2095.540 0.090 2103.340 2.700 ;
        RECT 2105.060 0.090 2112.860 2.700 ;
        RECT 2114.580 0.090 2122.380 2.700 ;
        RECT 2124.100 0.090 2131.900 2.700 ;
        RECT 2133.620 0.090 2141.420 2.700 ;
        RECT 2143.140 0.090 2150.940 2.700 ;
        RECT 2152.660 0.090 2160.460 2.700 ;
        RECT 2162.180 0.090 2169.980 2.700 ;
        RECT 2171.700 0.090 2179.500 2.700 ;
        RECT 2181.220 0.090 2189.020 2.700 ;
        RECT 2190.740 0.090 2198.540 2.700 ;
        RECT 2200.260 0.090 2208.060 2.700 ;
        RECT 2209.780 0.090 2217.580 2.700 ;
        RECT 2219.300 0.090 2227.100 2.700 ;
        RECT 2228.820 0.090 2236.620 2.700 ;
        RECT 2238.340 0.090 2246.140 2.700 ;
        RECT 2247.860 0.090 2255.660 2.700 ;
        RECT 2257.380 0.090 2265.180 2.700 ;
        RECT 2266.900 0.090 2274.700 2.700 ;
        RECT 2276.420 0.090 2284.220 2.700 ;
        RECT 2285.940 0.090 2293.740 2.700 ;
        RECT 2295.460 0.090 2303.260 2.700 ;
        RECT 2304.980 0.090 2312.780 2.700 ;
        RECT 2314.500 0.090 2322.300 2.700 ;
        RECT 2324.020 0.090 2331.820 2.700 ;
        RECT 2333.540 0.090 2341.340 2.700 ;
        RECT 2343.060 0.090 2350.860 2.700 ;
        RECT 2352.580 0.090 2360.380 2.700 ;
        RECT 2362.100 0.090 2369.900 2.700 ;
        RECT 2371.620 0.090 2379.420 2.700 ;
        RECT 2381.140 0.090 2388.940 2.700 ;
        RECT 2390.660 0.090 2398.460 2.700 ;
        RECT 2400.180 0.090 2407.980 2.700 ;
        RECT 2409.700 0.090 2417.500 2.700 ;
        RECT 2419.220 0.090 2427.020 2.700 ;
        RECT 2428.740 0.090 2436.540 2.700 ;
        RECT 2438.260 0.090 2446.060 2.700 ;
        RECT 2447.780 0.090 2455.580 2.700 ;
        RECT 2457.300 0.090 2465.100 2.700 ;
        RECT 2466.820 0.090 2474.620 2.700 ;
        RECT 2476.340 0.090 2484.140 2.700 ;
        RECT 2485.860 0.090 2493.660 2.700 ;
        RECT 2495.380 0.090 2503.180 2.700 ;
        RECT 2504.900 0.090 2512.700 2.700 ;
        RECT 2514.420 0.090 2522.220 2.700 ;
        RECT 2523.940 0.090 2531.740 2.700 ;
        RECT 2533.460 0.090 2541.260 2.700 ;
        RECT 2542.980 0.090 2550.780 2.700 ;
        RECT 2552.500 0.090 2560.300 2.700 ;
        RECT 2562.020 0.090 2569.820 2.700 ;
        RECT 2571.540 0.090 2579.340 2.700 ;
        RECT 2581.060 0.090 2588.860 2.700 ;
        RECT 2590.580 0.090 2598.380 2.700 ;
        RECT 2600.100 0.090 2607.900 2.700 ;
        RECT 2609.620 0.090 2617.420 2.700 ;
        RECT 2619.140 0.090 2626.940 2.700 ;
        RECT 2628.660 0.090 2636.460 2.700 ;
        RECT 2638.180 0.090 2645.980 2.700 ;
        RECT 2647.700 0.090 2655.500 2.700 ;
        RECT 2657.220 0.090 2665.020 2.700 ;
        RECT 2666.740 0.090 2674.540 2.700 ;
        RECT 2676.260 0.090 2684.060 2.700 ;
        RECT 2685.780 0.090 2693.580 2.700 ;
        RECT 2695.300 0.090 2703.100 2.700 ;
        RECT 2704.820 0.090 2712.620 2.700 ;
        RECT 2714.340 0.090 2722.140 2.700 ;
        RECT 2723.860 0.090 2731.660 2.700 ;
        RECT 2733.380 0.090 2741.180 2.700 ;
        RECT 2742.900 0.090 2750.700 2.700 ;
        RECT 2752.420 0.090 2760.220 2.700 ;
        RECT 2761.940 0.090 2769.740 2.700 ;
        RECT 2771.460 0.090 2779.260 2.700 ;
        RECT 2780.980 0.090 2788.780 2.700 ;
        RECT 2790.500 0.090 2798.300 2.700 ;
        RECT 2800.020 0.090 2807.820 2.700 ;
        RECT 2809.540 0.090 2817.340 2.700 ;
        RECT 2819.060 0.090 2826.860 2.700 ;
        RECT 2828.580 0.090 2836.380 2.700 ;
        RECT 2838.100 0.090 2845.900 2.700 ;
        RECT 2847.620 0.090 2855.420 2.700 ;
        RECT 2857.140 0.090 2864.940 2.700 ;
        RECT 2866.660 0.090 2874.460 2.700 ;
        RECT 2876.180 0.090 2883.980 2.700 ;
        RECT 2885.700 0.090 2893.500 2.700 ;
        RECT 2895.220 0.090 2903.020 2.700 ;
        RECT 2904.740 0.090 2912.540 2.700 ;
        RECT 2914.260 0.090 2922.060 2.700 ;
        RECT 2923.780 0.090 2931.580 2.700 ;
        RECT 2933.300 0.090 2992.500 2.700 ;
      LAYER Metal3 ;
        RECT 1.820 2966.900 2998.100 2979.060 ;
        RECT 1.820 2965.180 2997.300 2966.900 ;
        RECT 1.820 2958.500 2998.100 2965.180 ;
        RECT 2.700 2956.780 2998.100 2958.500 ;
        RECT 1.820 2900.260 2998.100 2956.780 ;
        RECT 1.820 2898.540 2997.300 2900.260 ;
        RECT 1.820 2887.380 2998.100 2898.540 ;
        RECT 2.700 2885.660 2998.100 2887.380 ;
        RECT 1.820 2833.620 2998.100 2885.660 ;
        RECT 1.820 2831.900 2997.300 2833.620 ;
        RECT 1.820 2816.260 2998.100 2831.900 ;
        RECT 2.700 2814.540 2998.100 2816.260 ;
        RECT 1.820 2766.980 2998.100 2814.540 ;
        RECT 1.820 2765.260 2997.300 2766.980 ;
        RECT 1.820 2745.140 2998.100 2765.260 ;
        RECT 2.700 2743.420 2998.100 2745.140 ;
        RECT 1.820 2700.340 2998.100 2743.420 ;
        RECT 1.820 2698.620 2997.300 2700.340 ;
        RECT 1.820 2674.020 2998.100 2698.620 ;
        RECT 2.700 2672.300 2998.100 2674.020 ;
        RECT 1.820 2633.700 2998.100 2672.300 ;
        RECT 1.820 2631.980 2997.300 2633.700 ;
        RECT 1.820 2602.900 2998.100 2631.980 ;
        RECT 2.700 2601.180 2998.100 2602.900 ;
        RECT 1.820 2567.060 2998.100 2601.180 ;
        RECT 1.820 2565.340 2997.300 2567.060 ;
        RECT 1.820 2531.780 2998.100 2565.340 ;
        RECT 2.700 2530.060 2998.100 2531.780 ;
        RECT 1.820 2500.420 2998.100 2530.060 ;
        RECT 1.820 2498.700 2997.300 2500.420 ;
        RECT 1.820 2460.660 2998.100 2498.700 ;
        RECT 2.700 2458.940 2998.100 2460.660 ;
        RECT 1.820 2433.780 2998.100 2458.940 ;
        RECT 1.820 2432.060 2997.300 2433.780 ;
        RECT 1.820 2389.540 2998.100 2432.060 ;
        RECT 2.700 2387.820 2998.100 2389.540 ;
        RECT 1.820 2367.140 2998.100 2387.820 ;
        RECT 1.820 2365.420 2997.300 2367.140 ;
        RECT 1.820 2318.420 2998.100 2365.420 ;
        RECT 2.700 2316.700 2998.100 2318.420 ;
        RECT 1.820 2300.500 2998.100 2316.700 ;
        RECT 1.820 2298.780 2997.300 2300.500 ;
        RECT 1.820 2247.300 2998.100 2298.780 ;
        RECT 2.700 2245.580 2998.100 2247.300 ;
        RECT 1.820 2233.860 2998.100 2245.580 ;
        RECT 1.820 2232.140 2997.300 2233.860 ;
        RECT 1.820 2176.180 2998.100 2232.140 ;
        RECT 2.700 2174.460 2998.100 2176.180 ;
        RECT 1.820 2167.220 2998.100 2174.460 ;
        RECT 1.820 2165.500 2997.300 2167.220 ;
        RECT 1.820 2105.060 2998.100 2165.500 ;
        RECT 2.700 2103.340 2998.100 2105.060 ;
        RECT 1.820 2100.580 2998.100 2103.340 ;
        RECT 1.820 2098.860 2997.300 2100.580 ;
        RECT 1.820 2033.940 2998.100 2098.860 ;
        RECT 2.700 2032.220 2997.300 2033.940 ;
        RECT 1.820 1967.300 2998.100 2032.220 ;
        RECT 1.820 1965.580 2997.300 1967.300 ;
        RECT 1.820 1962.820 2998.100 1965.580 ;
        RECT 2.700 1961.100 2998.100 1962.820 ;
        RECT 1.820 1900.660 2998.100 1961.100 ;
        RECT 1.820 1898.940 2997.300 1900.660 ;
        RECT 1.820 1891.700 2998.100 1898.940 ;
        RECT 2.700 1889.980 2998.100 1891.700 ;
        RECT 1.820 1834.020 2998.100 1889.980 ;
        RECT 1.820 1832.300 2997.300 1834.020 ;
        RECT 1.820 1820.580 2998.100 1832.300 ;
        RECT 2.700 1818.860 2998.100 1820.580 ;
        RECT 1.820 1767.380 2998.100 1818.860 ;
        RECT 1.820 1765.660 2997.300 1767.380 ;
        RECT 1.820 1749.460 2998.100 1765.660 ;
        RECT 2.700 1747.740 2998.100 1749.460 ;
        RECT 1.820 1700.740 2998.100 1747.740 ;
        RECT 1.820 1699.020 2997.300 1700.740 ;
        RECT 1.820 1678.340 2998.100 1699.020 ;
        RECT 2.700 1676.620 2998.100 1678.340 ;
        RECT 1.820 1634.100 2998.100 1676.620 ;
        RECT 1.820 1632.380 2997.300 1634.100 ;
        RECT 1.820 1607.220 2998.100 1632.380 ;
        RECT 2.700 1605.500 2998.100 1607.220 ;
        RECT 1.820 1567.460 2998.100 1605.500 ;
        RECT 1.820 1565.740 2997.300 1567.460 ;
        RECT 1.820 1536.100 2998.100 1565.740 ;
        RECT 2.700 1534.380 2998.100 1536.100 ;
        RECT 1.820 1500.820 2998.100 1534.380 ;
        RECT 1.820 1499.100 2997.300 1500.820 ;
        RECT 1.820 1464.980 2998.100 1499.100 ;
        RECT 2.700 1463.260 2998.100 1464.980 ;
        RECT 1.820 1434.180 2998.100 1463.260 ;
        RECT 1.820 1432.460 2997.300 1434.180 ;
        RECT 1.820 1393.860 2998.100 1432.460 ;
        RECT 2.700 1392.140 2998.100 1393.860 ;
        RECT 1.820 1367.540 2998.100 1392.140 ;
        RECT 1.820 1365.820 2997.300 1367.540 ;
        RECT 1.820 1322.740 2998.100 1365.820 ;
        RECT 2.700 1321.020 2998.100 1322.740 ;
        RECT 1.820 1300.900 2998.100 1321.020 ;
        RECT 1.820 1299.180 2997.300 1300.900 ;
        RECT 1.820 1251.620 2998.100 1299.180 ;
        RECT 2.700 1249.900 2998.100 1251.620 ;
        RECT 1.820 1234.260 2998.100 1249.900 ;
        RECT 1.820 1232.540 2997.300 1234.260 ;
        RECT 1.820 1180.500 2998.100 1232.540 ;
        RECT 2.700 1178.780 2998.100 1180.500 ;
        RECT 1.820 1167.620 2998.100 1178.780 ;
        RECT 1.820 1165.900 2997.300 1167.620 ;
        RECT 1.820 1109.380 2998.100 1165.900 ;
        RECT 2.700 1107.660 2998.100 1109.380 ;
        RECT 1.820 1100.980 2998.100 1107.660 ;
        RECT 1.820 1099.260 2997.300 1100.980 ;
        RECT 1.820 1038.260 2998.100 1099.260 ;
        RECT 2.700 1036.540 2998.100 1038.260 ;
        RECT 1.820 1034.340 2998.100 1036.540 ;
        RECT 1.820 1032.620 2997.300 1034.340 ;
        RECT 1.820 967.700 2998.100 1032.620 ;
        RECT 1.820 967.140 2997.300 967.700 ;
        RECT 2.700 965.980 2997.300 967.140 ;
        RECT 2.700 965.420 2998.100 965.980 ;
        RECT 1.820 901.060 2998.100 965.420 ;
        RECT 1.820 899.340 2997.300 901.060 ;
        RECT 1.820 896.020 2998.100 899.340 ;
        RECT 2.700 894.300 2998.100 896.020 ;
        RECT 1.820 834.420 2998.100 894.300 ;
        RECT 1.820 832.700 2997.300 834.420 ;
        RECT 1.820 824.900 2998.100 832.700 ;
        RECT 2.700 823.180 2998.100 824.900 ;
        RECT 1.820 767.780 2998.100 823.180 ;
        RECT 1.820 766.060 2997.300 767.780 ;
        RECT 1.820 753.780 2998.100 766.060 ;
        RECT 2.700 752.060 2998.100 753.780 ;
        RECT 1.820 701.140 2998.100 752.060 ;
        RECT 1.820 699.420 2997.300 701.140 ;
        RECT 1.820 682.660 2998.100 699.420 ;
        RECT 2.700 680.940 2998.100 682.660 ;
        RECT 1.820 634.500 2998.100 680.940 ;
        RECT 1.820 632.780 2997.300 634.500 ;
        RECT 1.820 611.540 2998.100 632.780 ;
        RECT 2.700 609.820 2998.100 611.540 ;
        RECT 1.820 567.860 2998.100 609.820 ;
        RECT 1.820 566.140 2997.300 567.860 ;
        RECT 1.820 540.420 2998.100 566.140 ;
        RECT 2.700 538.700 2998.100 540.420 ;
        RECT 1.820 501.220 2998.100 538.700 ;
        RECT 1.820 499.500 2997.300 501.220 ;
        RECT 1.820 469.300 2998.100 499.500 ;
        RECT 2.700 467.580 2998.100 469.300 ;
        RECT 1.820 434.580 2998.100 467.580 ;
        RECT 1.820 432.860 2997.300 434.580 ;
        RECT 1.820 398.180 2998.100 432.860 ;
        RECT 2.700 396.460 2998.100 398.180 ;
        RECT 1.820 367.940 2998.100 396.460 ;
        RECT 1.820 366.220 2997.300 367.940 ;
        RECT 1.820 327.060 2998.100 366.220 ;
        RECT 2.700 325.340 2998.100 327.060 ;
        RECT 1.820 301.300 2998.100 325.340 ;
        RECT 1.820 299.580 2997.300 301.300 ;
        RECT 1.820 255.940 2998.100 299.580 ;
        RECT 2.700 254.220 2998.100 255.940 ;
        RECT 1.820 234.660 2998.100 254.220 ;
        RECT 1.820 232.940 2997.300 234.660 ;
        RECT 1.820 184.820 2998.100 232.940 ;
        RECT 2.700 183.100 2998.100 184.820 ;
        RECT 1.820 168.020 2998.100 183.100 ;
        RECT 1.820 166.300 2997.300 168.020 ;
        RECT 1.820 113.700 2998.100 166.300 ;
        RECT 2.700 111.980 2998.100 113.700 ;
        RECT 1.820 101.380 2998.100 111.980 ;
        RECT 1.820 99.660 2997.300 101.380 ;
        RECT 1.820 42.580 2998.100 99.660 ;
        RECT 2.700 40.860 2998.100 42.580 ;
        RECT 1.820 34.740 2998.100 40.860 ;
        RECT 1.820 33.020 2997.300 34.740 ;
        RECT 1.820 0.140 2998.100 33.020 ;
      LAYER Metal4 ;
        RECT 398.860 20.250 403.590 2978.550 ;
        RECT 407.290 20.250 474.990 2978.550 ;
        RECT 478.690 20.250 493.590 2978.550 ;
        RECT 497.290 20.250 564.990 2978.550 ;
        RECT 568.690 20.250 583.590 2978.550 ;
        RECT 587.290 20.250 654.990 2978.550 ;
        RECT 658.690 20.250 673.590 2978.550 ;
        RECT 677.290 20.250 744.990 2978.550 ;
        RECT 748.690 20.250 763.590 2978.550 ;
        RECT 767.290 20.250 834.990 2978.550 ;
        RECT 838.690 20.250 853.590 2978.550 ;
        RECT 857.290 20.250 924.990 2978.550 ;
        RECT 928.690 20.250 943.590 2978.550 ;
        RECT 947.290 20.250 1014.990 2978.550 ;
        RECT 1018.690 1344.280 1033.590 2978.550 ;
        RECT 1037.290 1344.280 1104.990 2978.550 ;
        RECT 1018.690 555.400 1104.990 1344.280 ;
        RECT 1018.690 20.250 1033.590 555.400 ;
        RECT 1037.290 20.250 1104.990 555.400 ;
        RECT 1108.690 20.250 1123.590 2978.550 ;
        RECT 1127.290 20.250 1194.990 2978.550 ;
        RECT 1198.690 20.250 1213.590 2978.550 ;
        RECT 1217.290 20.250 1284.990 2978.550 ;
        RECT 1288.690 20.250 1303.590 2978.550 ;
        RECT 1307.290 20.250 1374.990 2978.550 ;
        RECT 1378.690 20.250 1393.590 2978.550 ;
        RECT 1397.290 20.250 1464.990 2978.550 ;
        RECT 1468.690 20.250 1483.590 2978.550 ;
        RECT 1487.290 20.250 1501.220 2978.550 ;
  END
END user_project_wrapper
END LIBRARY

